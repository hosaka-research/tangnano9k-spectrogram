module nco_rom (clock,ce,oce,reset,addr,dataout);
	input clock,ce,oce,reset;
	input [8:0] addr;
	output [17:0] dataout;
	reg [17:0] dataout;
	always @(posedge clock or posedge reset) begin
		if(reset) begin
			dataout <= 0;
		end else begin
			if (ce & oce) begin
				case (addr)
					9'h0000: dataout<=18'h1ece6;
					9'h0001: dataout<=18'h08a86;
					9'h0002: dataout<=18'h1fb33;
					9'h0003: dataout<=18'h045ea;
					9'h0004: dataout<=18'h1ea94;
					9'h0005: dataout<=18'h09289;
					9'h0006: dataout<=18'h1fa9d;
					9'h0007: dataout<=18'h04a0b;
					9'h0008: dataout<=18'h1e7f9;
					9'h0009: dataout<=18'h09afb;
					9'h000a: dataout<=18'h1f9f4;
					9'h000b: dataout<=18'h04e6a;
					9'h000c: dataout<=18'h00000;
					9'h000d: dataout<=18'h00000;
					9'h000e: dataout<=18'h00000;
					9'h000f: dataout<=18'h00000;
					9'h0010: dataout<=18'h00000;
					9'h0011: dataout<=18'h00000;
					9'h0012: dataout<=18'h00000;
					9'h0013: dataout<=18'h00000;
					9'h0014: dataout<=18'h00000;
					9'h0015: dataout<=18'h00000;
					9'h0016: dataout<=18'h00000;
					9'h0017: dataout<=18'h00000;
					9'h0018: dataout<=18'h00000;
					9'h0019: dataout<=18'h00000;
					9'h001a: dataout<=18'h00000;
					9'h001b: dataout<=18'h00000;
					9'h001c: dataout<=18'h00000;
					9'h001d: dataout<=18'h00000;
					9'h001e: dataout<=18'h00000;
					9'h001f: dataout<=18'h00000;
					9'h0020: dataout<=18'h00000;
					9'h0021: dataout<=18'h00000;
					9'h0022: dataout<=18'h00000;
					9'h0023: dataout<=18'h00000;
					9'h0024: dataout<=18'h00000;
					9'h0025: dataout<=18'h00000;
					9'h0026: dataout<=18'h00000;
					9'h0027: dataout<=18'h00000;
					9'h0028: dataout<=18'h00000;
					9'h0029: dataout<=18'h00000;
					9'h002a: dataout<=18'h00000;
					9'h002b: dataout<=18'h00000;
					9'h002c: dataout<=18'h00000;
					9'h002d: dataout<=18'h00000;
					9'h002e: dataout<=18'h00000;
					9'h002f: dataout<=18'h00000;
					9'h0030: dataout<=18'h00000;
					9'h0031: dataout<=18'h00000;
					9'h0032: dataout<=18'h00000;
					9'h0033: dataout<=18'h00000;
					9'h0034: dataout<=18'h00000;
					9'h0035: dataout<=18'h00000;
					9'h0036: dataout<=18'h00000;
					9'h0037: dataout<=18'h00000;
					9'h0038: dataout<=18'h00000;
					9'h0039: dataout<=18'h00000;
					9'h003a: dataout<=18'h00000;
					9'h003b: dataout<=18'h00000;
					9'h003c: dataout<=18'h00000;
					9'h003d: dataout<=18'h00000;
					9'h003e: dataout<=18'h00000;
					9'h003f: dataout<=18'h00000;
					9'h0040: dataout<=18'h00000;
					9'h0041: dataout<=18'h00000;
					9'h0042: dataout<=18'h00000;
					9'h0043: dataout<=18'h00000;
					9'h0044: dataout<=18'h00000;
					9'h0045: dataout<=18'h00000;
					9'h0046: dataout<=18'h00000;
					9'h0047: dataout<=18'h00000;
					9'h0048: dataout<=18'h00000;
					9'h0049: dataout<=18'h00000;
					9'h004a: dataout<=18'h00000;
					9'h004b: dataout<=18'h00000;
					9'h004c: dataout<=18'h00000;
					9'h004d: dataout<=18'h00000;
					9'h004e: dataout<=18'h00000;
					9'h004f: dataout<=18'h00000;
					9'h0050: dataout<=18'h00000;
					9'h0051: dataout<=18'h00000;
					9'h0052: dataout<=18'h00000;
					9'h0053: dataout<=18'h00000;
					9'h0054: dataout<=18'h00000;
					9'h0055: dataout<=18'h00000;
					9'h0056: dataout<=18'h00000;
					9'h0057: dataout<=18'h00000;
					9'h0058: dataout<=18'h00000;
					9'h0059: dataout<=18'h00000;
					9'h005a: dataout<=18'h00000;
					9'h005b: dataout<=18'h00000;
					9'h005c: dataout<=18'h00000;
					9'h005d: dataout<=18'h00000;
					9'h005e: dataout<=18'h00000;
					9'h005f: dataout<=18'h00000;
					9'h0060: dataout<=18'h00000;
					9'h0061: dataout<=18'h00000;
					9'h0062: dataout<=18'h00000;
					9'h0063: dataout<=18'h00000;
					9'h0064: dataout<=18'h00000;
					9'h0065: dataout<=18'h00000;
					9'h0066: dataout<=18'h00000;
					9'h0067: dataout<=18'h00000;
					9'h0068: dataout<=18'h00000;
					9'h0069: dataout<=18'h00000;
					9'h006a: dataout<=18'h00000;
					9'h006b: dataout<=18'h00000;
					9'h006c: dataout<=18'h00000;
					9'h006d: dataout<=18'h00000;
					9'h006e: dataout<=18'h00000;
					9'h006f: dataout<=18'h00000;
					9'h0070: dataout<=18'h00000;
					9'h0071: dataout<=18'h00000;
					9'h0072: dataout<=18'h00000;
					9'h0073: dataout<=18'h00000;
					9'h0074: dataout<=18'h00000;
					9'h0075: dataout<=18'h00000;
					9'h0076: dataout<=18'h00000;
					9'h0077: dataout<=18'h00000;
					9'h0078: dataout<=18'h00000;
					9'h0079: dataout<=18'h00000;
					9'h007a: dataout<=18'h00000;
					9'h007b: dataout<=18'h00000;
					9'h007c: dataout<=18'h00000;
					9'h007d: dataout<=18'h00000;
					9'h007e: dataout<=18'h00000;
					9'h007f: dataout<=18'h00000;
					9'h0080: dataout<=18'h00000;
					9'h0081: dataout<=18'h00000;
					9'h0082: dataout<=18'h00000;
					9'h0083: dataout<=18'h00000;
					9'h0084: dataout<=18'h00000;
					9'h0085: dataout<=18'h00000;
					9'h0086: dataout<=18'h00000;
					9'h0087: dataout<=18'h00000;
					9'h0088: dataout<=18'h00000;
					9'h0089: dataout<=18'h00000;
					9'h008a: dataout<=18'h00000;
					9'h008b: dataout<=18'h00000;
					9'h008c: dataout<=18'h00000;
					9'h008d: dataout<=18'h00000;
					9'h008e: dataout<=18'h00000;
					9'h008f: dataout<=18'h00000;
					9'h0090: dataout<=18'h00000;
					9'h0091: dataout<=18'h00000;
					9'h0092: dataout<=18'h00000;
					9'h0093: dataout<=18'h00000;
					9'h0094: dataout<=18'h00000;
					9'h0095: dataout<=18'h00000;
					9'h0096: dataout<=18'h00000;
					9'h0097: dataout<=18'h00000;
					9'h0098: dataout<=18'h00000;
					9'h0099: dataout<=18'h00000;
					9'h009a: dataout<=18'h00000;
					9'h009b: dataout<=18'h00000;
					9'h009c: dataout<=18'h00000;
					9'h009d: dataout<=18'h00000;
					9'h009e: dataout<=18'h00000;
					9'h009f: dataout<=18'h00000;
					9'h00a0: dataout<=18'h00000;
					9'h00a1: dataout<=18'h00000;
					9'h00a2: dataout<=18'h00000;
					9'h00a3: dataout<=18'h00000;
					9'h00a4: dataout<=18'h00000;
					9'h00a5: dataout<=18'h00000;
					9'h00a6: dataout<=18'h00000;
					9'h00a7: dataout<=18'h00000;
					9'h00a8: dataout<=18'h00000;
					9'h00a9: dataout<=18'h00000;
					9'h00aa: dataout<=18'h00000;
					9'h00ab: dataout<=18'h00000;
					9'h00ac: dataout<=18'h00000;
					9'h00ad: dataout<=18'h00000;
					9'h00ae: dataout<=18'h00000;
					9'h00af: dataout<=18'h00000;
					9'h00b0: dataout<=18'h00000;
					9'h00b1: dataout<=18'h00000;
					9'h00b2: dataout<=18'h00000;
					9'h00b3: dataout<=18'h00000;
					9'h00b4: dataout<=18'h00000;
					9'h00b5: dataout<=18'h00000;
					9'h00b6: dataout<=18'h00000;
					9'h00b7: dataout<=18'h00000;
					9'h00b8: dataout<=18'h00000;
					9'h00b9: dataout<=18'h00000;
					9'h00ba: dataout<=18'h00000;
					9'h00bb: dataout<=18'h00000;
					9'h00bc: dataout<=18'h00000;
					9'h00bd: dataout<=18'h00000;
					9'h00be: dataout<=18'h00000;
					9'h00bf: dataout<=18'h00000;
					9'h00c0: dataout<=18'h00000;
					9'h00c1: dataout<=18'h00000;
					9'h00c2: dataout<=18'h00000;
					9'h00c3: dataout<=18'h00000;
					9'h00c4: dataout<=18'h00000;
					9'h00c5: dataout<=18'h00000;
					9'h00c6: dataout<=18'h00000;
					9'h00c7: dataout<=18'h00000;
					9'h00c8: dataout<=18'h00000;
					9'h00c9: dataout<=18'h00000;
					9'h00ca: dataout<=18'h00000;
					9'h00cb: dataout<=18'h00000;
					9'h00cc: dataout<=18'h00000;
					9'h00cd: dataout<=18'h00000;
					9'h00ce: dataout<=18'h00000;
					9'h00cf: dataout<=18'h00000;
					9'h00d0: dataout<=18'h00000;
					9'h00d1: dataout<=18'h00000;
					9'h00d2: dataout<=18'h00000;
					9'h00d3: dataout<=18'h00000;
					9'h00d4: dataout<=18'h00000;
					9'h00d5: dataout<=18'h00000;
					9'h00d6: dataout<=18'h00000;
					9'h00d7: dataout<=18'h00000;
					9'h00d8: dataout<=18'h00000;
					9'h00d9: dataout<=18'h00000;
					9'h00da: dataout<=18'h00000;
					9'h00db: dataout<=18'h00000;
					9'h00dc: dataout<=18'h00000;
					9'h00dd: dataout<=18'h00000;
					9'h00de: dataout<=18'h00000;
					9'h00df: dataout<=18'h00000;
					9'h00e0: dataout<=18'h00000;
					9'h00e1: dataout<=18'h00000;
					9'h00e2: dataout<=18'h00000;
					9'h00e3: dataout<=18'h00000;
					9'h00e4: dataout<=18'h00000;
					9'h00e5: dataout<=18'h00000;
					9'h00e6: dataout<=18'h00000;
					9'h00e7: dataout<=18'h00000;
					9'h00e8: dataout<=18'h00000;
					9'h00e9: dataout<=18'h00000;
					9'h00ea: dataout<=18'h00000;
					9'h00eb: dataout<=18'h00000;
					9'h00ec: dataout<=18'h00000;
					9'h00ed: dataout<=18'h00000;
					9'h00ee: dataout<=18'h00000;
					9'h00ef: dataout<=18'h00000;
					9'h00f0: dataout<=18'h00000;
					9'h00f1: dataout<=18'h00000;
					9'h00f2: dataout<=18'h00000;
					9'h00f3: dataout<=18'h00000;
					9'h00f4: dataout<=18'h00000;
					9'h00f5: dataout<=18'h00000;
					9'h00f6: dataout<=18'h00000;
					9'h00f7: dataout<=18'h00000;
					9'h00f8: dataout<=18'h00000;
					9'h00f9: dataout<=18'h00000;
					9'h00fa: dataout<=18'h00000;
					9'h00fb: dataout<=18'h00000;
					9'h00fc: dataout<=18'h00000;
					9'h00fd: dataout<=18'h00000;
					9'h00fe: dataout<=18'h00000;
					9'h00ff: dataout<=18'h00000;
					9'h0100: dataout<=18'h00000;
					9'h0101: dataout<=18'h00000;
					9'h0102: dataout<=18'h00000;
					9'h0103: dataout<=18'h00000;
					9'h0104: dataout<=18'h00000;
					9'h0105: dataout<=18'h00000;
					9'h0106: dataout<=18'h00000;
					9'h0107: dataout<=18'h00000;
					9'h0108: dataout<=18'h00000;
					9'h0109: dataout<=18'h00000;
					9'h010a: dataout<=18'h00000;
					9'h010b: dataout<=18'h00000;
					9'h010c: dataout<=18'h00000;
					9'h010d: dataout<=18'h00000;
					9'h010e: dataout<=18'h00000;
					9'h010f: dataout<=18'h00000;
					9'h0110: dataout<=18'h00000;
					9'h0111: dataout<=18'h00000;
					9'h0112: dataout<=18'h00000;
					9'h0113: dataout<=18'h00000;
					9'h0114: dataout<=18'h00000;
					9'h0115: dataout<=18'h00000;
					9'h0116: dataout<=18'h00000;
					9'h0117: dataout<=18'h00000;
					9'h0118: dataout<=18'h00000;
					9'h0119: dataout<=18'h00000;
					9'h011a: dataout<=18'h00000;
					9'h011b: dataout<=18'h00000;
					9'h011c: dataout<=18'h00000;
					9'h011d: dataout<=18'h00000;
					9'h011e: dataout<=18'h00000;
					9'h011f: dataout<=18'h00000;
					9'h0120: dataout<=18'h00000;
					9'h0121: dataout<=18'h00000;
					9'h0122: dataout<=18'h00000;
					9'h0123: dataout<=18'h00000;
					9'h0124: dataout<=18'h00000;
					9'h0125: dataout<=18'h00000;
					9'h0126: dataout<=18'h00000;
					9'h0127: dataout<=18'h00000;
					9'h0128: dataout<=18'h00000;
					9'h0129: dataout<=18'h00000;
					9'h012a: dataout<=18'h00000;
					9'h012b: dataout<=18'h00000;
					9'h012c: dataout<=18'h00000;
					9'h012d: dataout<=18'h00000;
					9'h012e: dataout<=18'h00000;
					9'h012f: dataout<=18'h00000;
					9'h0130: dataout<=18'h00000;
					9'h0131: dataout<=18'h00000;
					9'h0132: dataout<=18'h00000;
					9'h0133: dataout<=18'h00000;
					9'h0134: dataout<=18'h00000;
					9'h0135: dataout<=18'h00000;
					9'h0136: dataout<=18'h00000;
					9'h0137: dataout<=18'h00000;
					9'h0138: dataout<=18'h00000;
					9'h0139: dataout<=18'h00000;
					9'h013a: dataout<=18'h00000;
					9'h013b: dataout<=18'h00000;
					9'h013c: dataout<=18'h00000;
					9'h013d: dataout<=18'h00000;
					9'h013e: dataout<=18'h00000;
					9'h013f: dataout<=18'h00000;
					9'h0140: dataout<=18'h00000;
					9'h0141: dataout<=18'h00000;
					9'h0142: dataout<=18'h00000;
					9'h0143: dataout<=18'h00000;
					9'h0144: dataout<=18'h00000;
					9'h0145: dataout<=18'h00000;
					9'h0146: dataout<=18'h00000;
					9'h0147: dataout<=18'h00000;
					9'h0148: dataout<=18'h00000;
					9'h0149: dataout<=18'h00000;
					9'h014a: dataout<=18'h00000;
					9'h014b: dataout<=18'h00000;
					9'h014c: dataout<=18'h00000;
					9'h014d: dataout<=18'h00000;
					9'h014e: dataout<=18'h00000;
					9'h014f: dataout<=18'h00000;
					9'h0150: dataout<=18'h00000;
					9'h0151: dataout<=18'h00000;
					9'h0152: dataout<=18'h00000;
					9'h0153: dataout<=18'h00000;
					9'h0154: dataout<=18'h00000;
					9'h0155: dataout<=18'h00000;
					9'h0156: dataout<=18'h00000;
					9'h0157: dataout<=18'h00000;
					9'h0158: dataout<=18'h00000;
					9'h0159: dataout<=18'h00000;
					9'h015a: dataout<=18'h00000;
					9'h015b: dataout<=18'h00000;
					9'h015c: dataout<=18'h00000;
					9'h015d: dataout<=18'h00000;
					9'h015e: dataout<=18'h00000;
					9'h015f: dataout<=18'h00000;
					9'h0160: dataout<=18'h00000;
					9'h0161: dataout<=18'h00000;
					9'h0162: dataout<=18'h00000;
					9'h0163: dataout<=18'h00000;
					9'h0164: dataout<=18'h00000;
					9'h0165: dataout<=18'h00000;
					9'h0166: dataout<=18'h00000;
					9'h0167: dataout<=18'h00000;
					9'h0168: dataout<=18'h00000;
					9'h0169: dataout<=18'h00000;
					9'h016a: dataout<=18'h00000;
					9'h016b: dataout<=18'h00000;
					9'h016c: dataout<=18'h00000;
					9'h016d: dataout<=18'h00000;
					9'h016e: dataout<=18'h00000;
					9'h016f: dataout<=18'h00000;
					9'h0170: dataout<=18'h00000;
					9'h0171: dataout<=18'h00000;
					9'h0172: dataout<=18'h00000;
					9'h0173: dataout<=18'h00000;
					9'h0174: dataout<=18'h00000;
					9'h0175: dataout<=18'h00000;
					9'h0176: dataout<=18'h00000;
					9'h0177: dataout<=18'h00000;
					9'h0178: dataout<=18'h00000;
					9'h0179: dataout<=18'h00000;
					9'h017a: dataout<=18'h00000;
					9'h017b: dataout<=18'h00000;
					9'h017c: dataout<=18'h00000;
					9'h017d: dataout<=18'h00000;
					9'h017e: dataout<=18'h00000;
					9'h017f: dataout<=18'h00000;
					9'h0180: dataout<=18'h00000;
					9'h0181: dataout<=18'h00000;
					9'h0182: dataout<=18'h00000;
					9'h0183: dataout<=18'h00000;
					9'h0184: dataout<=18'h00000;
					9'h0185: dataout<=18'h00000;
					9'h0186: dataout<=18'h00000;
					9'h0187: dataout<=18'h00000;
					9'h0188: dataout<=18'h00000;
					9'h0189: dataout<=18'h00000;
					9'h018a: dataout<=18'h00000;
					9'h018b: dataout<=18'h00000;
					9'h018c: dataout<=18'h00000;
					9'h018d: dataout<=18'h00000;
					9'h018e: dataout<=18'h00000;
					9'h018f: dataout<=18'h00000;
					9'h0190: dataout<=18'h00000;
					9'h0191: dataout<=18'h00000;
					9'h0192: dataout<=18'h00000;
					9'h0193: dataout<=18'h00000;
					9'h0194: dataout<=18'h00000;
					9'h0195: dataout<=18'h00000;
					9'h0196: dataout<=18'h00000;
					9'h0197: dataout<=18'h00000;
					9'h0198: dataout<=18'h00000;
					9'h0199: dataout<=18'h00000;
					9'h019a: dataout<=18'h00000;
					9'h019b: dataout<=18'h00000;
					9'h019c: dataout<=18'h00000;
					9'h019d: dataout<=18'h00000;
					9'h019e: dataout<=18'h00000;
					9'h019f: dataout<=18'h00000;
					9'h01a0: dataout<=18'h00000;
					9'h01a1: dataout<=18'h00000;
					9'h01a2: dataout<=18'h00000;
					9'h01a3: dataout<=18'h00000;
					9'h01a4: dataout<=18'h00000;
					9'h01a5: dataout<=18'h00000;
					9'h01a6: dataout<=18'h00000;
					9'h01a7: dataout<=18'h00000;
					9'h01a8: dataout<=18'h00000;
					9'h01a9: dataout<=18'h00000;
					9'h01aa: dataout<=18'h00000;
					9'h01ab: dataout<=18'h00000;
					9'h01ac: dataout<=18'h00000;
					9'h01ad: dataout<=18'h00000;
					9'h01ae: dataout<=18'h00000;
					9'h01af: dataout<=18'h00000;
					9'h01b0: dataout<=18'h00000;
					9'h01b1: dataout<=18'h00000;
					9'h01b2: dataout<=18'h00000;
					9'h01b3: dataout<=18'h00000;
					9'h01b4: dataout<=18'h00000;
					9'h01b5: dataout<=18'h00000;
					9'h01b6: dataout<=18'h00000;
					9'h01b7: dataout<=18'h00000;
					9'h01b8: dataout<=18'h00000;
					9'h01b9: dataout<=18'h00000;
					9'h01ba: dataout<=18'h00000;
					9'h01bb: dataout<=18'h00000;
					9'h01bc: dataout<=18'h00000;
					9'h01bd: dataout<=18'h00000;
					9'h01be: dataout<=18'h00000;
					9'h01bf: dataout<=18'h00000;
					9'h01c0: dataout<=18'h00000;
					9'h01c1: dataout<=18'h00000;
					9'h01c2: dataout<=18'h00000;
					9'h01c3: dataout<=18'h00000;
					9'h01c4: dataout<=18'h00000;
					9'h01c5: dataout<=18'h00000;
					9'h01c6: dataout<=18'h00000;
					9'h01c7: dataout<=18'h00000;
					9'h01c8: dataout<=18'h00000;
					9'h01c9: dataout<=18'h00000;
					9'h01ca: dataout<=18'h00000;
					9'h01cb: dataout<=18'h00000;
					9'h01cc: dataout<=18'h00000;
					9'h01cd: dataout<=18'h00000;
					9'h01ce: dataout<=18'h00000;
					9'h01cf: dataout<=18'h00000;
					9'h01d0: dataout<=18'h00000;
					9'h01d1: dataout<=18'h00000;
					9'h01d2: dataout<=18'h00000;
					9'h01d3: dataout<=18'h00000;
					9'h01d4: dataout<=18'h00000;
					9'h01d5: dataout<=18'h00000;
					9'h01d6: dataout<=18'h00000;
					9'h01d7: dataout<=18'h00000;
					9'h01d8: dataout<=18'h00000;
					9'h01d9: dataout<=18'h00000;
					9'h01da: dataout<=18'h00000;
					9'h01db: dataout<=18'h00000;
					9'h01dc: dataout<=18'h00000;
					9'h01dd: dataout<=18'h00000;
					9'h01de: dataout<=18'h00000;
					9'h01df: dataout<=18'h00000;
					9'h01e0: dataout<=18'h00000;
					9'h01e1: dataout<=18'h00000;
					9'h01e2: dataout<=18'h00000;
					9'h01e3: dataout<=18'h00000;
					9'h01e4: dataout<=18'h00000;
					9'h01e5: dataout<=18'h00000;
					9'h01e6: dataout<=18'h00000;
					9'h01e7: dataout<=18'h00000;
					9'h01e8: dataout<=18'h00000;
					9'h01e9: dataout<=18'h00000;
					9'h01ea: dataout<=18'h00000;
					9'h01eb: dataout<=18'h00000;
					9'h01ec: dataout<=18'h00000;
					9'h01ed: dataout<=18'h00000;
					9'h01ee: dataout<=18'h00000;
					9'h01ef: dataout<=18'h00000;
					9'h01f0: dataout<=18'h00000;
					9'h01f1: dataout<=18'h00000;
					9'h01f2: dataout<=18'h00000;
					9'h01f3: dataout<=18'h00000;
					9'h01f4: dataout<=18'h00000;
					9'h01f5: dataout<=18'h00000;
					9'h01f6: dataout<=18'h00000;
					9'h01f7: dataout<=18'h00000;
					9'h01f8: dataout<=18'h00000;
					9'h01f9: dataout<=18'h00000;
					9'h01fa: dataout<=18'h00000;
					9'h01fb: dataout<=18'h00000;
					9'h01fc: dataout<=18'h00000;
					9'h01fd: dataout<=18'h00000;
					9'h01fe: dataout<=18'h00000;
					9'h01ff: dataout<=18'h00000;
				endcase
			end
		end
	end
endmodule

