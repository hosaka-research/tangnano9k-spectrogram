module fctheta_rom (clock,ce,oce,reset,addr,dataout);
	input clock,ce,oce,reset;
	input [9:0] addr;
	output [35:0] dataout;
	reg [35:0] dataout;
	always @(posedge clock or posedge reset) begin
		if(reset) begin
			dataout <= 0;
		end else begin
			if (ce & oce) begin
				case (addr)
					10'd0000: dataout<=36'd27487790694;
					10'd0001: dataout<=36'd27430644017;
					10'd0002: dataout<=36'd27373497340;
					10'd0003: dataout<=36'd27316350663;
					10'd0004: dataout<=36'd27259203986;
					10'd0005: dataout<=36'd27202057309;
					10'd0006: dataout<=36'd27144910633;
					10'd0007: dataout<=36'd27087763956;
					10'd0008: dataout<=36'd27030617279;
					10'd0009: dataout<=36'd26973470602;
					10'd0010: dataout<=36'd26916323925;
					10'd0011: dataout<=36'd26859177248;
					10'd0012: dataout<=36'd26802030571;
					10'd0013: dataout<=36'd26744883894;
					10'd0014: dataout<=36'd26687737217;
					10'd0015: dataout<=36'd26630590540;
					10'd0016: dataout<=36'd26573443864;
					10'd0017: dataout<=36'd26516297187;
					10'd0018: dataout<=36'd26459150510;
					10'd0019: dataout<=36'd26402003833;
					10'd0020: dataout<=36'd26344857156;
					10'd0021: dataout<=36'd26287710479;
					10'd0022: dataout<=36'd26230563802;
					10'd0023: dataout<=36'd26173417125;
					10'd0024: dataout<=36'd26116270448;
					10'd0025: dataout<=36'd26059123772;
					10'd0026: dataout<=36'd26001977095;
					10'd0027: dataout<=36'd25944830418;
					10'd0028: dataout<=36'd25887683741;
					10'd0029: dataout<=36'd25830537064;
					10'd0030: dataout<=36'd25773390387;
					10'd0031: dataout<=36'd25716243710;
					10'd0032: dataout<=36'd25659097033;
					10'd0033: dataout<=36'd25601950356;
					10'd0034: dataout<=36'd25544803679;
					10'd0035: dataout<=36'd25487657003;
					10'd0036: dataout<=36'd25430510326;
					10'd0037: dataout<=36'd25373363649;
					10'd0038: dataout<=36'd25316216972;
					10'd0039: dataout<=36'd25259070295;
					10'd0040: dataout<=36'd25201923618;
					10'd0041: dataout<=36'd25144776941;
					10'd0042: dataout<=36'd25087630264;
					10'd0043: dataout<=36'd25030483587;
					10'd0044: dataout<=36'd24973336910;
					10'd0045: dataout<=36'd24916190234;
					10'd0046: dataout<=36'd24859043557;
					10'd0047: dataout<=36'd24801896880;
					10'd0048: dataout<=36'd24744750203;
					10'd0049: dataout<=36'd24687603526;
					10'd0050: dataout<=36'd24630456849;
					10'd0051: dataout<=36'd24573310172;
					10'd0052: dataout<=36'd24516163495;
					10'd0053: dataout<=36'd24459016818;
					10'd0054: dataout<=36'd24401870142;
					10'd0055: dataout<=36'd24344723465;
					10'd0056: dataout<=36'd24287576788;
					10'd0057: dataout<=36'd24230430111;
					10'd0058: dataout<=36'd24173283434;
					10'd0059: dataout<=36'd24116136757;
					10'd0060: dataout<=36'd24058990080;
					10'd0061: dataout<=36'd24001843403;
					10'd0062: dataout<=36'd23944696726;
					10'd0063: dataout<=36'd23887550049;
					10'd0064: dataout<=36'd23830403373;
					10'd0065: dataout<=36'd23773256696;
					10'd0066: dataout<=36'd23716110019;
					10'd0067: dataout<=36'd23658963342;
					10'd0068: dataout<=36'd23601816665;
					10'd0069: dataout<=36'd23544669988;
					10'd0070: dataout<=36'd23487523311;
					10'd0071: dataout<=36'd23430376634;
					10'd0072: dataout<=36'd23373229957;
					10'd0073: dataout<=36'd23316083280;
					10'd0074: dataout<=36'd23258936604;
					10'd0075: dataout<=36'd23201789927;
					10'd0076: dataout<=36'd23144643250;
					10'd0077: dataout<=36'd23087496573;
					10'd0078: dataout<=36'd23030349896;
					10'd0079: dataout<=36'd22973203219;
					10'd0080: dataout<=36'd22916056542;
					10'd0081: dataout<=36'd22858909865;
					10'd0082: dataout<=36'd22801763188;
					10'd0083: dataout<=36'd22744616512;
					10'd0084: dataout<=36'd22687469835;
					10'd0085: dataout<=36'd22630323158;
					10'd0086: dataout<=36'd22573176481;
					10'd0087: dataout<=36'd22516029804;
					10'd0088: dataout<=36'd22458883127;
					10'd0089: dataout<=36'd22401736450;
					10'd0090: dataout<=36'd22344589773;
					10'd0091: dataout<=36'd22287443096;
					10'd0092: dataout<=36'd22230296419;
					10'd0093: dataout<=36'd22173149743;
					10'd0094: dataout<=36'd22116003066;
					10'd0095: dataout<=36'd22058856389;
					10'd0096: dataout<=36'd22001709712;
					10'd0097: dataout<=36'd21944563035;
					10'd0098: dataout<=36'd21887416358;
					10'd0099: dataout<=36'd21830269681;
					10'd0100: dataout<=36'd21773123004;
					10'd0101: dataout<=36'd21715976327;
					10'd0102: dataout<=36'd21658829651;
					10'd0103: dataout<=36'd21601682974;
					10'd0104: dataout<=36'd21544536297;
					10'd0105: dataout<=36'd21487389620;
					10'd0106: dataout<=36'd21430242943;
					10'd0107: dataout<=36'd21373096266;
					10'd0108: dataout<=36'd21315949589;
					10'd0109: dataout<=36'd21258802912;
					10'd0110: dataout<=36'd21201656235;
					10'd0111: dataout<=36'd21144509558;
					10'd0112: dataout<=36'd21087362882;
					10'd0113: dataout<=36'd21030216205;
					10'd0114: dataout<=36'd20973069528;
					10'd0115: dataout<=36'd20915922851;
					10'd0116: dataout<=36'd20858776174;
					10'd0117: dataout<=36'd20801629497;
					10'd0118: dataout<=36'd20744482820;
					10'd0119: dataout<=36'd20687336143;
					10'd0120: dataout<=36'd20630189466;
					10'd0121: dataout<=36'd20573042789;
					10'd0122: dataout<=36'd20515896113;
					10'd0123: dataout<=36'd20458749436;
					10'd0124: dataout<=36'd20401602759;
					10'd0125: dataout<=36'd20344456082;
					10'd0126: dataout<=36'd20287309405;
					10'd0127: dataout<=36'd20230162728;
					10'd0128: dataout<=36'd20173016051;
					10'd0129: dataout<=36'd20115869374;
					10'd0130: dataout<=36'd20058722697;
					10'd0131: dataout<=36'd20001576021;
					10'd0132: dataout<=36'd19944429344;
					10'd0133: dataout<=36'd19887282667;
					10'd0134: dataout<=36'd19830135990;
					10'd0135: dataout<=36'd19772989313;
					10'd0136: dataout<=36'd19715842636;
					10'd0137: dataout<=36'd19658695959;
					10'd0138: dataout<=36'd19601549282;
					10'd0139: dataout<=36'd19544402605;
					10'd0140: dataout<=36'd19487255928;
					10'd0141: dataout<=36'd19430109252;
					10'd0142: dataout<=36'd19372962575;
					10'd0143: dataout<=36'd19315815898;
					10'd0144: dataout<=36'd19258669221;
					10'd0145: dataout<=36'd19201522544;
					10'd0146: dataout<=36'd19144375867;
					10'd0147: dataout<=36'd19087229190;
					10'd0148: dataout<=36'd19030082513;
					10'd0149: dataout<=36'd18972935836;
					10'd0150: dataout<=36'd18915789160;
					10'd0151: dataout<=36'd18858642483;
					10'd0152: dataout<=36'd18801495806;
					10'd0153: dataout<=36'd18744349129;
					10'd0154: dataout<=36'd18687202452;
					10'd0155: dataout<=36'd18630055775;
					10'd0156: dataout<=36'd18572909098;
					10'd0157: dataout<=36'd18515762421;
					10'd0158: dataout<=36'd18458615744;
					10'd0159: dataout<=36'd18401469067;
					10'd0160: dataout<=36'd18344322391;
					10'd0161: dataout<=36'd18287175714;
					10'd0162: dataout<=36'd18230029037;
					10'd0163: dataout<=36'd18172882360;
					10'd0164: dataout<=36'd18115735683;
					10'd0165: dataout<=36'd18058589006;
					10'd0166: dataout<=36'd18001442329;
					10'd0167: dataout<=36'd17944295652;
					10'd0168: dataout<=36'd17887148975;
					10'd0169: dataout<=36'd17830002298;
					10'd0170: dataout<=36'd17772855622;
					10'd0171: dataout<=36'd17715708945;
					10'd0172: dataout<=36'd17658562268;
					10'd0173: dataout<=36'd17601415591;
					10'd0174: dataout<=36'd17544268914;
					10'd0175: dataout<=36'd17487122237;
					10'd0176: dataout<=36'd17429975560;
					10'd0177: dataout<=36'd17372828883;
					10'd0178: dataout<=36'd17315682206;
					10'd0179: dataout<=36'd17258535530;
					10'd0180: dataout<=36'd17201388853;
					10'd0181: dataout<=36'd17144242176;
					10'd0182: dataout<=36'd17087095499;
					10'd0183: dataout<=36'd17029948822;
					10'd0184: dataout<=36'd16972802145;
					10'd0185: dataout<=36'd16915655468;
					10'd0186: dataout<=36'd16858508791;
					10'd0187: dataout<=36'd16801362114;
					10'd0188: dataout<=36'd16744215437;
					10'd0189: dataout<=36'd16687068761;
					10'd0190: dataout<=36'd16629922084;
					10'd0191: dataout<=36'd16572775407;
					10'd0192: dataout<=36'd16515628730;
					10'd0193: dataout<=36'd16458482053;
					10'd0194: dataout<=36'd16401335376;
					10'd0195: dataout<=36'd16344188699;
					10'd0196: dataout<=36'd16287042022;
					10'd0197: dataout<=36'd16229895345;
					10'd0198: dataout<=36'd16172748668;
					10'd0199: dataout<=36'd16115601992;
					10'd0200: dataout<=36'd16058455315;
					10'd0201: dataout<=36'd16001308638;
					10'd0202: dataout<=36'd15944161961;
					10'd0203: dataout<=36'd15887015284;
					10'd0204: dataout<=36'd15829868607;
					10'd0205: dataout<=36'd15772721930;
					10'd0206: dataout<=36'd15715575253;
					10'd0207: dataout<=36'd15658428576;
					10'd0208: dataout<=36'd15601281900;
					10'd0209: dataout<=36'd15544135223;
					10'd0210: dataout<=36'd15486988546;
					10'd0211: dataout<=36'd15429841869;
					10'd0212: dataout<=36'd15372695192;
					10'd0213: dataout<=36'd15315548515;
					10'd0214: dataout<=36'd15258401838;
					10'd0215: dataout<=36'd15201255161;
					10'd0216: dataout<=36'd15144108484;
					10'd0217: dataout<=36'd15086961807;
					10'd0218: dataout<=36'd15029815131;
					10'd0219: dataout<=36'd14972668454;
					10'd0220: dataout<=36'd14915521777;
					10'd0221: dataout<=36'd14858375100;
					10'd0222: dataout<=36'd14801228423;
					10'd0223: dataout<=36'd14744081746;
					10'd0224: dataout<=36'd14686935069;
					10'd0225: dataout<=36'd14629788392;
					10'd0226: dataout<=36'd14572641715;
					10'd0227: dataout<=36'd14515495039;
					10'd0228: dataout<=36'd14458348362;
					10'd0229: dataout<=36'd14401201685;
					10'd0230: dataout<=36'd14344055008;
					10'd0231: dataout<=36'd14286908331;
					10'd0232: dataout<=36'd14229761654;
					10'd0233: dataout<=36'd14172614977;
					10'd0234: dataout<=36'd14115468300;
					10'd0235: dataout<=36'd14058321623;
					10'd0236: dataout<=36'd14001174946;
					10'd0237: dataout<=36'd13944028270;
					10'd0238: dataout<=36'd13886881593;
					10'd0239: dataout<=36'd13829734916;
					10'd0240: dataout<=36'd13772588239;
					10'd0241: dataout<=36'd13715441562;
					10'd0242: dataout<=36'd13658294885;
					10'd0243: dataout<=36'd13601148208;
					10'd0244: dataout<=36'd13544001531;
					10'd0245: dataout<=36'd13486854854;
					10'd0246: dataout<=36'd13429708177;
					10'd0247: dataout<=36'd13372561501;
					10'd0248: dataout<=36'd13315414824;
					10'd0249: dataout<=36'd13258268147;
					10'd0250: dataout<=36'd13201121470;
					10'd0251: dataout<=36'd13143974793;
					10'd0252: dataout<=36'd13086828116;
					10'd0253: dataout<=36'd13029681439;
					10'd0254: dataout<=36'd12972534762;
					10'd0255: dataout<=36'd12915388085;
					10'd0256: dataout<=36'd12858241409;
					10'd0257: dataout<=36'd12801094732;
					10'd0258: dataout<=36'd12743948055;
					10'd0259: dataout<=36'd12686801378;
					10'd0260: dataout<=36'd12629654701;
					10'd0261: dataout<=36'd12572508024;
					10'd0262: dataout<=36'd12515361347;
					10'd0263: dataout<=36'd12458214670;
					10'd0264: dataout<=36'd12401067993;
					10'd0265: dataout<=36'd12343921316;
					10'd0266: dataout<=36'd12286774640;
					10'd0267: dataout<=36'd12229627963;
					10'd0268: dataout<=36'd12172481286;
					10'd0269: dataout<=36'd12115334609;
					10'd0270: dataout<=36'd12058187932;
					10'd0271: dataout<=36'd12001041255;
					10'd0272: dataout<=36'd11943894578;
					10'd0273: dataout<=36'd11886747901;
					10'd0274: dataout<=36'd11829601224;
					10'd0275: dataout<=36'd11772454548;
					10'd0276: dataout<=36'd11715307871;
					10'd0277: dataout<=36'd11658161194;
					10'd0278: dataout<=36'd11601014517;
					10'd0279: dataout<=36'd11543867840;
					10'd0280: dataout<=36'd11486721163;
					10'd0281: dataout<=36'd11429574486;
					10'd0282: dataout<=36'd11372427809;
					10'd0283: dataout<=36'd11315281132;
					10'd0284: dataout<=36'd11258134455;
					10'd0285: dataout<=36'd11200987779;
					10'd0286: dataout<=36'd11143841102;
					10'd0287: dataout<=36'd11086694425;
					10'd0288: dataout<=36'd11029547748;
					10'd0289: dataout<=36'd10972401071;
					10'd0290: dataout<=36'd10915254394;
					10'd0291: dataout<=36'd10858107717;
					10'd0292: dataout<=36'd10800961040;
					10'd0293: dataout<=36'd10743814363;
					10'd0294: dataout<=36'd10686667686;
					10'd0295: dataout<=36'd10629521010;
					10'd0296: dataout<=36'd10572374333;
					10'd0297: dataout<=36'd10515227656;
					10'd0298: dataout<=36'd10458080979;
					10'd0299: dataout<=36'd10400934302;
					10'd0300: dataout<=36'd10343787625;
					10'd0301: dataout<=36'd10286640948;
					10'd0302: dataout<=36'd10229494271;
					10'd0303: dataout<=36'd10172347594;
					10'd0304: dataout<=36'd10115200918;
					10'd0305: dataout<=36'd10058054241;
					10'd0306: dataout<=36'd10000907564;
					10'd0307: dataout<=36'd9943760887;
					10'd0308: dataout<=36'd9886614210;
					10'd0309: dataout<=36'd9829467533;
					10'd0310: dataout<=36'd9772320856;
					10'd0311: dataout<=36'd9715174179;
					10'd0312: dataout<=36'd9658027502;
					10'd0313: dataout<=36'd9600880825;
					10'd0314: dataout<=36'd9543734149;
					10'd0315: dataout<=36'd9486587472;
					10'd0316: dataout<=36'd9429440795;
					10'd0317: dataout<=36'd9372294118;
					10'd0318: dataout<=36'd9315147441;
					10'd0319: dataout<=36'd9258000764;
					10'd0320: dataout<=36'd9200854087;
					10'd0321: dataout<=36'd9143707410;
					10'd0322: dataout<=36'd9086560733;
					10'd0323: dataout<=36'd9029414056;
					10'd0324: dataout<=36'd8972267380;
					10'd0325: dataout<=36'd8915120703;
					10'd0326: dataout<=36'd8857974026;
					10'd0327: dataout<=36'd8800827349;
					10'd0328: dataout<=36'd8743680672;
					10'd0329: dataout<=36'd8686533995;
					10'd0330: dataout<=36'd8629387318;
					10'd0331: dataout<=36'd8572240641;
					10'd0332: dataout<=36'd8515093964;
					10'd0333: dataout<=36'd8457947288;
					10'd0334: dataout<=36'd8400800611;
					10'd0335: dataout<=36'd8343653934;
					10'd0336: dataout<=36'd8286507257;
					10'd0337: dataout<=36'd8229360580;
					10'd0338: dataout<=36'd8172213903;
					10'd0339: dataout<=36'd8115067226;
					10'd0340: dataout<=36'd8057920549;
					10'd0341: dataout<=36'd8000773872;
					10'd0342: dataout<=36'd7943627195;
					10'd0343: dataout<=36'd7886480519;
					10'd0344: dataout<=36'd7829333842;
					10'd0345: dataout<=36'd7772187165;
					10'd0346: dataout<=36'd7715040488;
					10'd0347: dataout<=36'd7657893811;
					10'd0348: dataout<=36'd7600747134;
					10'd0349: dataout<=36'd7543600457;
					10'd0350: dataout<=36'd7486453780;
					10'd0351: dataout<=36'd7429307103;
					10'd0352: dataout<=36'd7372160427;
					10'd0353: dataout<=36'd7315013750;
					10'd0354: dataout<=36'd7257867073;
					10'd0355: dataout<=36'd7200720396;
					10'd0356: dataout<=36'd7143573719;
					10'd0357: dataout<=36'd7086427042;
					10'd0358: dataout<=36'd7029280365;
					10'd0359: dataout<=36'd6972133688;
					10'd0360: dataout<=36'd6914987011;
					10'd0361: dataout<=36'd6857840334;
					10'd0362: dataout<=36'd6800693658;
					10'd0363: dataout<=36'd6743546981;
					10'd0364: dataout<=36'd6686400304;
					10'd0365: dataout<=36'd6629253627;
					10'd0366: dataout<=36'd6572106950;
					10'd0367: dataout<=36'd6514960273;
					10'd0368: dataout<=36'd6457813596;
					10'd0369: dataout<=36'd6400666919;
					10'd0370: dataout<=36'd6343520242;
					10'd0371: dataout<=36'd6286373565;
					10'd0372: dataout<=36'd6229226889;
					10'd0373: dataout<=36'd6172080212;
					10'd0374: dataout<=36'd6114933535;
					10'd0375: dataout<=36'd6057786858;
					10'd0376: dataout<=36'd6000640181;
					10'd0377: dataout<=36'd5943493504;
					10'd0378: dataout<=36'd5886346827;
					10'd0379: dataout<=36'd5829200150;
					10'd0380: dataout<=36'd5772053473;
					10'd0381: dataout<=36'd5714906797;
					10'd0382: dataout<=36'd5657760120;
					10'd0383: dataout<=36'd5600613443;
					10'd0384: dataout<=36'd5543466766;
					10'd0385: dataout<=36'd5486320089;
					10'd0386: dataout<=36'd5429173412;
					10'd0387: dataout<=36'd5372026735;
					10'd0388: dataout<=36'd5314880058;
					10'd0389: dataout<=36'd5257733381;
					10'd0390: dataout<=36'd5200586704;
					10'd0391: dataout<=36'd5143440028;
					10'd0392: dataout<=36'd5086293351;
					10'd0393: dataout<=36'd5029146674;
					10'd0394: dataout<=36'd4971999997;
					10'd0395: dataout<=36'd4914853320;
					10'd0396: dataout<=36'd4857706643;
					10'd0397: dataout<=36'd4800559966;
					10'd0398: dataout<=36'd4743413289;
					10'd0399: dataout<=36'd4686266612;
					10'd0400: dataout<=36'd4629119936;
					10'd0401: dataout<=36'd4571973259;
					10'd0402: dataout<=36'd4514826582;
					10'd0403: dataout<=36'd4457679905;
					10'd0404: dataout<=36'd4400533228;
					10'd0405: dataout<=36'd4343386551;
					10'd0406: dataout<=36'd4286239874;
					10'd0407: dataout<=36'd4229093197;
					10'd0408: dataout<=36'd4171946520;
					10'd0409: dataout<=36'd4114799843;
					10'd0410: dataout<=36'd4057653167;
					10'd0411: dataout<=36'd4000506490;
					10'd0412: dataout<=36'd3943359813;
					10'd0413: dataout<=36'd3886213136;
					10'd0414: dataout<=36'd3829066459;
					10'd0415: dataout<=36'd3771919782;
					10'd0416: dataout<=36'd3714773105;
					10'd0417: dataout<=36'd3657626428;
					10'd0418: dataout<=36'd3600479751;
					10'd0419: dataout<=36'd3543333074;
					10'd0420: dataout<=36'd3486186398;
					10'd0421: dataout<=36'd3429039721;
					10'd0422: dataout<=36'd3371893044;
					10'd0423: dataout<=36'd3314746367;
					10'd0424: dataout<=36'd3257599690;
					10'd0425: dataout<=36'd3200453013;
					10'd0426: dataout<=36'd3143306336;
					10'd0427: dataout<=36'd3086159659;
					10'd0428: dataout<=36'd3029012982;
					10'd0429: dataout<=36'd2971866306;
					10'd0430: dataout<=36'd2914719629;
					10'd0431: dataout<=36'd2857572952;
					10'd0432: dataout<=36'd2800426275;
					10'd0433: dataout<=36'd2743279598;
					10'd0434: dataout<=36'd2686132921;
					10'd0435: dataout<=36'd2628986244;
					10'd0436: dataout<=36'd2571839567;
					10'd0437: dataout<=36'd2514692890;
					10'd0438: dataout<=36'd2457546213;
					10'd0439: dataout<=36'd2400399537;
					10'd0440: dataout<=36'd2343252860;
					10'd0441: dataout<=36'd2286106183;
					10'd0442: dataout<=36'd2228959506;
					10'd0443: dataout<=36'd2171812829;
					10'd0444: dataout<=36'd2114666152;
					10'd0445: dataout<=36'd2057519475;
					10'd0446: dataout<=36'd2000372798;
					10'd0447: dataout<=36'd1943226121;
					10'd0448: dataout<=36'd1886079445;
					10'd0449: dataout<=36'd1828932768;
					10'd0450: dataout<=36'd1771786091;
					10'd0451: dataout<=36'd1714639414;
					10'd0452: dataout<=36'd1657492737;
					10'd0453: dataout<=36'd1600346060;
					10'd0454: dataout<=36'd1543199383;
					10'd0455: dataout<=36'd1486052706;
					10'd0456: dataout<=36'd1428906029;
					10'd0457: dataout<=36'd1371759352;
					10'd0458: dataout<=36'd1314612676;
					10'd0459: dataout<=36'd1257465999;
					10'd0460: dataout<=36'd1200319322;
					10'd0461: dataout<=36'd1143172645;
					10'd0462: dataout<=36'd1086025968;
					10'd0463: dataout<=36'd1028879291;
					10'd0464: dataout<=36'd971732614;
					10'd0465: dataout<=36'd914585937;
					10'd0466: dataout<=36'd857439260;
					10'd0467: dataout<=36'd800292583;
					10'd0468: dataout<=36'd743145907;
					10'd0469: dataout<=36'd685999230;
					10'd0470: dataout<=36'd628852553;
					10'd0471: dataout<=36'd571705876;
					10'd0472: dataout<=36'd514559199;
					10'd0473: dataout<=36'd457412522;
					10'd0474: dataout<=36'd400265845;
					10'd0475: dataout<=36'd343119168;
					10'd0476: dataout<=36'd285972491;
					10'd0477: dataout<=36'd228825815;
					10'd0478: dataout<=36'd171679138;
					10'd0479: dataout<=36'd114532461;
					10'd0480: dataout<=36'd00000000;
					10'd0481: dataout<=36'd00000000;
					10'd0482: dataout<=36'd00000000;
					10'd0483: dataout<=36'd00000000;
					10'd0484: dataout<=36'd00000000;
					10'd0485: dataout<=36'd00000000;
					10'd0486: dataout<=36'd00000000;
					10'd0487: dataout<=36'd00000000;
					10'd0488: dataout<=36'd00000000;
					10'd0489: dataout<=36'd00000000;
					10'd0490: dataout<=36'd00000000;
					10'd0491: dataout<=36'd00000000;
					10'd0492: dataout<=36'd00000000;
					10'd0493: dataout<=36'd00000000;
					10'd0494: dataout<=36'd00000000;
					10'd0495: dataout<=36'd00000000;
					10'd0496: dataout<=36'd00000000;
					10'd0497: dataout<=36'd00000000;
					10'd0498: dataout<=36'd00000000;
					10'd0499: dataout<=36'd00000000;
					10'd0500: dataout<=36'd00000000;
					10'd0501: dataout<=36'd00000000;
					10'd0502: dataout<=36'd00000000;
					10'd0503: dataout<=36'd00000000;
					10'd0504: dataout<=36'd00000000;
					10'd0505: dataout<=36'd00000000;
					10'd0506: dataout<=36'd00000000;
					10'd0507: dataout<=36'd00000000;
					10'd0508: dataout<=36'd00000000;
					10'd0509: dataout<=36'd00000000;
					10'd0510: dataout<=36'd00000000;
					10'd0511: dataout<=36'd00000000;
					10'd0512: dataout<=36'd00000000;
					10'd0513: dataout<=36'd00000000;
					10'd0514: dataout<=36'd00000000;
					10'd0515: dataout<=36'd00000000;
					10'd0516: dataout<=36'd00000000;
					10'd0517: dataout<=36'd00000000;
					10'd0518: dataout<=36'd00000000;
					10'd0519: dataout<=36'd00000000;
					10'd0520: dataout<=36'd00000000;
					10'd0521: dataout<=36'd00000000;
					10'd0522: dataout<=36'd00000000;
					10'd0523: dataout<=36'd00000000;
					10'd0524: dataout<=36'd00000000;
					10'd0525: dataout<=36'd00000000;
					10'd0526: dataout<=36'd00000000;
					10'd0527: dataout<=36'd00000000;
					10'd0528: dataout<=36'd00000000;
					10'd0529: dataout<=36'd00000000;
					10'd0530: dataout<=36'd00000000;
					10'd0531: dataout<=36'd00000000;
					10'd0532: dataout<=36'd00000000;
					10'd0533: dataout<=36'd00000000;
					10'd0534: dataout<=36'd00000000;
					10'd0535: dataout<=36'd00000000;
					10'd0536: dataout<=36'd00000000;
					10'd0537: dataout<=36'd00000000;
					10'd0538: dataout<=36'd00000000;
					10'd0539: dataout<=36'd00000000;
					10'd0540: dataout<=36'd00000000;
					10'd0541: dataout<=36'd00000000;
					10'd0542: dataout<=36'd00000000;
					10'd0543: dataout<=36'd00000000;
					10'd0544: dataout<=36'd00000000;
					10'd0545: dataout<=36'd00000000;
					10'd0546: dataout<=36'd00000000;
					10'd0547: dataout<=36'd00000000;
					10'd0548: dataout<=36'd00000000;
					10'd0549: dataout<=36'd00000000;
					10'd0550: dataout<=36'd00000000;
					10'd0551: dataout<=36'd00000000;
					10'd0552: dataout<=36'd00000000;
					10'd0553: dataout<=36'd00000000;
					10'd0554: dataout<=36'd00000000;
					10'd0555: dataout<=36'd00000000;
					10'd0556: dataout<=36'd00000000;
					10'd0557: dataout<=36'd00000000;
					10'd0558: dataout<=36'd00000000;
					10'd0559: dataout<=36'd00000000;
					10'd0560: dataout<=36'd00000000;
					10'd0561: dataout<=36'd00000000;
					10'd0562: dataout<=36'd00000000;
					10'd0563: dataout<=36'd00000000;
					10'd0564: dataout<=36'd00000000;
					10'd0565: dataout<=36'd00000000;
					10'd0566: dataout<=36'd00000000;
					10'd0567: dataout<=36'd00000000;
					10'd0568: dataout<=36'd00000000;
					10'd0569: dataout<=36'd00000000;
					10'd0570: dataout<=36'd00000000;
					10'd0571: dataout<=36'd00000000;
					10'd0572: dataout<=36'd00000000;
					10'd0573: dataout<=36'd00000000;
					10'd0574: dataout<=36'd00000000;
					10'd0575: dataout<=36'd00000000;
					10'd0576: dataout<=36'd00000000;
					10'd0577: dataout<=36'd00000000;
					10'd0578: dataout<=36'd00000000;
					10'd0579: dataout<=36'd00000000;
					10'd0580: dataout<=36'd00000000;
					10'd0581: dataout<=36'd00000000;
					10'd0582: dataout<=36'd00000000;
					10'd0583: dataout<=36'd00000000;
					10'd0584: dataout<=36'd00000000;
					10'd0585: dataout<=36'd00000000;
					10'd0586: dataout<=36'd00000000;
					10'd0587: dataout<=36'd00000000;
					10'd0588: dataout<=36'd00000000;
					10'd0589: dataout<=36'd00000000;
					10'd0590: dataout<=36'd00000000;
					10'd0591: dataout<=36'd00000000;
					10'd0592: dataout<=36'd00000000;
					10'd0593: dataout<=36'd00000000;
					10'd0594: dataout<=36'd00000000;
					10'd0595: dataout<=36'd00000000;
					10'd0596: dataout<=36'd00000000;
					10'd0597: dataout<=36'd00000000;
					10'd0598: dataout<=36'd00000000;
					10'd0599: dataout<=36'd00000000;
					10'd0600: dataout<=36'd00000000;
					10'd0601: dataout<=36'd00000000;
					10'd0602: dataout<=36'd00000000;
					10'd0603: dataout<=36'd00000000;
					10'd0604: dataout<=36'd00000000;
					10'd0605: dataout<=36'd00000000;
					10'd0606: dataout<=36'd00000000;
					10'd0607: dataout<=36'd00000000;
					10'd0608: dataout<=36'd00000000;
					10'd0609: dataout<=36'd00000000;
					10'd0610: dataout<=36'd00000000;
					10'd0611: dataout<=36'd00000000;
					10'd0612: dataout<=36'd00000000;
					10'd0613: dataout<=36'd00000000;
					10'd0614: dataout<=36'd00000000;
					10'd0615: dataout<=36'd00000000;
					10'd0616: dataout<=36'd00000000;
					10'd0617: dataout<=36'd00000000;
					10'd0618: dataout<=36'd00000000;
					10'd0619: dataout<=36'd00000000;
					10'd0620: dataout<=36'd00000000;
					10'd0621: dataout<=36'd00000000;
					10'd0622: dataout<=36'd00000000;
					10'd0623: dataout<=36'd00000000;
					10'd0624: dataout<=36'd00000000;
					10'd0625: dataout<=36'd00000000;
					10'd0626: dataout<=36'd00000000;
					10'd0627: dataout<=36'd00000000;
					10'd0628: dataout<=36'd00000000;
					10'd0629: dataout<=36'd00000000;
					10'd0630: dataout<=36'd00000000;
					10'd0631: dataout<=36'd00000000;
					10'd0632: dataout<=36'd00000000;
					10'd0633: dataout<=36'd00000000;
					10'd0634: dataout<=36'd00000000;
					10'd0635: dataout<=36'd00000000;
					10'd0636: dataout<=36'd00000000;
					10'd0637: dataout<=36'd00000000;
					10'd0638: dataout<=36'd00000000;
					10'd0639: dataout<=36'd00000000;
					10'd0640: dataout<=36'd00000000;
					10'd0641: dataout<=36'd00000000;
					10'd0642: dataout<=36'd00000000;
					10'd0643: dataout<=36'd00000000;
					10'd0644: dataout<=36'd00000000;
					10'd0645: dataout<=36'd00000000;
					10'd0646: dataout<=36'd00000000;
					10'd0647: dataout<=36'd00000000;
					10'd0648: dataout<=36'd00000000;
					10'd0649: dataout<=36'd00000000;
					10'd0650: dataout<=36'd00000000;
					10'd0651: dataout<=36'd00000000;
					10'd0652: dataout<=36'd00000000;
					10'd0653: dataout<=36'd00000000;
					10'd0654: dataout<=36'd00000000;
					10'd0655: dataout<=36'd00000000;
					10'd0656: dataout<=36'd00000000;
					10'd0657: dataout<=36'd00000000;
					10'd0658: dataout<=36'd00000000;
					10'd0659: dataout<=36'd00000000;
					10'd0660: dataout<=36'd00000000;
					10'd0661: dataout<=36'd00000000;
					10'd0662: dataout<=36'd00000000;
					10'd0663: dataout<=36'd00000000;
					10'd0664: dataout<=36'd00000000;
					10'd0665: dataout<=36'd00000000;
					10'd0666: dataout<=36'd00000000;
					10'd0667: dataout<=36'd00000000;
					10'd0668: dataout<=36'd00000000;
					10'd0669: dataout<=36'd00000000;
					10'd0670: dataout<=36'd00000000;
					10'd0671: dataout<=36'd00000000;
					10'd0672: dataout<=36'd00000000;
					10'd0673: dataout<=36'd00000000;
					10'd0674: dataout<=36'd00000000;
					10'd0675: dataout<=36'd00000000;
					10'd0676: dataout<=36'd00000000;
					10'd0677: dataout<=36'd00000000;
					10'd0678: dataout<=36'd00000000;
					10'd0679: dataout<=36'd00000000;
					10'd0680: dataout<=36'd00000000;
					10'd0681: dataout<=36'd00000000;
					10'd0682: dataout<=36'd00000000;
					10'd0683: dataout<=36'd00000000;
					10'd0684: dataout<=36'd00000000;
					10'd0685: dataout<=36'd00000000;
					10'd0686: dataout<=36'd00000000;
					10'd0687: dataout<=36'd00000000;
					10'd0688: dataout<=36'd00000000;
					10'd0689: dataout<=36'd00000000;
					10'd0690: dataout<=36'd00000000;
					10'd0691: dataout<=36'd00000000;
					10'd0692: dataout<=36'd00000000;
					10'd0693: dataout<=36'd00000000;
					10'd0694: dataout<=36'd00000000;
					10'd0695: dataout<=36'd00000000;
					10'd0696: dataout<=36'd00000000;
					10'd0697: dataout<=36'd00000000;
					10'd0698: dataout<=36'd00000000;
					10'd0699: dataout<=36'd00000000;
					10'd0700: dataout<=36'd00000000;
					10'd0701: dataout<=36'd00000000;
					10'd0702: dataout<=36'd00000000;
					10'd0703: dataout<=36'd00000000;
					10'd0704: dataout<=36'd00000000;
					10'd0705: dataout<=36'd00000000;
					10'd0706: dataout<=36'd00000000;
					10'd0707: dataout<=36'd00000000;
					10'd0708: dataout<=36'd00000000;
					10'd0709: dataout<=36'd00000000;
					10'd0710: dataout<=36'd00000000;
					10'd0711: dataout<=36'd00000000;
					10'd0712: dataout<=36'd00000000;
					10'd0713: dataout<=36'd00000000;
					10'd0714: dataout<=36'd00000000;
					10'd0715: dataout<=36'd00000000;
					10'd0716: dataout<=36'd00000000;
					10'd0717: dataout<=36'd00000000;
					10'd0718: dataout<=36'd00000000;
					10'd0719: dataout<=36'd00000000;
					10'd0720: dataout<=36'd00000000;
					10'd0721: dataout<=36'd00000000;
					10'd0722: dataout<=36'd00000000;
					10'd0723: dataout<=36'd00000000;
					10'd0724: dataout<=36'd00000000;
					10'd0725: dataout<=36'd00000000;
					10'd0726: dataout<=36'd00000000;
					10'd0727: dataout<=36'd00000000;
					10'd0728: dataout<=36'd00000000;
					10'd0729: dataout<=36'd00000000;
					10'd0730: dataout<=36'd00000000;
					10'd0731: dataout<=36'd00000000;
					10'd0732: dataout<=36'd00000000;
					10'd0733: dataout<=36'd00000000;
					10'd0734: dataout<=36'd00000000;
					10'd0735: dataout<=36'd00000000;
					10'd0736: dataout<=36'd00000000;
					10'd0737: dataout<=36'd00000000;
					10'd0738: dataout<=36'd00000000;
					10'd0739: dataout<=36'd00000000;
					10'd0740: dataout<=36'd00000000;
					10'd0741: dataout<=36'd00000000;
					10'd0742: dataout<=36'd00000000;
					10'd0743: dataout<=36'd00000000;
					10'd0744: dataout<=36'd00000000;
					10'd0745: dataout<=36'd00000000;
					10'd0746: dataout<=36'd00000000;
					10'd0747: dataout<=36'd00000000;
					10'd0748: dataout<=36'd00000000;
					10'd0749: dataout<=36'd00000000;
					10'd0750: dataout<=36'd00000000;
					10'd0751: dataout<=36'd00000000;
					10'd0752: dataout<=36'd00000000;
					10'd0753: dataout<=36'd00000000;
					10'd0754: dataout<=36'd00000000;
					10'd0755: dataout<=36'd00000000;
					10'd0756: dataout<=36'd00000000;
					10'd0757: dataout<=36'd00000000;
					10'd0758: dataout<=36'd00000000;
					10'd0759: dataout<=36'd00000000;
					10'd0760: dataout<=36'd00000000;
					10'd0761: dataout<=36'd00000000;
					10'd0762: dataout<=36'd00000000;
					10'd0763: dataout<=36'd00000000;
					10'd0764: dataout<=36'd00000000;
					10'd0765: dataout<=36'd00000000;
					10'd0766: dataout<=36'd00000000;
					10'd0767: dataout<=36'd00000000;
					10'd0768: dataout<=36'd00000000;
					10'd0769: dataout<=36'd00000000;
					10'd0770: dataout<=36'd00000000;
					10'd0771: dataout<=36'd00000000;
					10'd0772: dataout<=36'd00000000;
					10'd0773: dataout<=36'd00000000;
					10'd0774: dataout<=36'd00000000;
					10'd0775: dataout<=36'd00000000;
					10'd0776: dataout<=36'd00000000;
					10'd0777: dataout<=36'd00000000;
					10'd0778: dataout<=36'd00000000;
					10'd0779: dataout<=36'd00000000;
					10'd0780: dataout<=36'd00000000;
					10'd0781: dataout<=36'd00000000;
					10'd0782: dataout<=36'd00000000;
					10'd0783: dataout<=36'd00000000;
					10'd0784: dataout<=36'd00000000;
					10'd0785: dataout<=36'd00000000;
					10'd0786: dataout<=36'd00000000;
					10'd0787: dataout<=36'd00000000;
					10'd0788: dataout<=36'd00000000;
					10'd0789: dataout<=36'd00000000;
					10'd0790: dataout<=36'd00000000;
					10'd0791: dataout<=36'd00000000;
					10'd0792: dataout<=36'd00000000;
					10'd0793: dataout<=36'd00000000;
					10'd0794: dataout<=36'd00000000;
					10'd0795: dataout<=36'd00000000;
					10'd0796: dataout<=36'd00000000;
					10'd0797: dataout<=36'd00000000;
					10'd0798: dataout<=36'd00000000;
					10'd0799: dataout<=36'd00000000;
					10'd0800: dataout<=36'd00000000;
					10'd0801: dataout<=36'd00000000;
					10'd0802: dataout<=36'd00000000;
					10'd0803: dataout<=36'd00000000;
					10'd0804: dataout<=36'd00000000;
					10'd0805: dataout<=36'd00000000;
					10'd0806: dataout<=36'd00000000;
					10'd0807: dataout<=36'd00000000;
					10'd0808: dataout<=36'd00000000;
					10'd0809: dataout<=36'd00000000;
					10'd0810: dataout<=36'd00000000;
					10'd0811: dataout<=36'd00000000;
					10'd0812: dataout<=36'd00000000;
					10'd0813: dataout<=36'd00000000;
					10'd0814: dataout<=36'd00000000;
					10'd0815: dataout<=36'd00000000;
					10'd0816: dataout<=36'd00000000;
					10'd0817: dataout<=36'd00000000;
					10'd0818: dataout<=36'd00000000;
					10'd0819: dataout<=36'd00000000;
					10'd0820: dataout<=36'd00000000;
					10'd0821: dataout<=36'd00000000;
					10'd0822: dataout<=36'd00000000;
					10'd0823: dataout<=36'd00000000;
					10'd0824: dataout<=36'd00000000;
					10'd0825: dataout<=36'd00000000;
					10'd0826: dataout<=36'd00000000;
					10'd0827: dataout<=36'd00000000;
					10'd0828: dataout<=36'd00000000;
					10'd0829: dataout<=36'd00000000;
					10'd0830: dataout<=36'd00000000;
					10'd0831: dataout<=36'd00000000;
					10'd0832: dataout<=36'd00000000;
					10'd0833: dataout<=36'd00000000;
					10'd0834: dataout<=36'd00000000;
					10'd0835: dataout<=36'd00000000;
					10'd0836: dataout<=36'd00000000;
					10'd0837: dataout<=36'd00000000;
					10'd0838: dataout<=36'd00000000;
					10'd0839: dataout<=36'd00000000;
					10'd0840: dataout<=36'd00000000;
					10'd0841: dataout<=36'd00000000;
					10'd0842: dataout<=36'd00000000;
					10'd0843: dataout<=36'd00000000;
					10'd0844: dataout<=36'd00000000;
					10'd0845: dataout<=36'd00000000;
					10'd0846: dataout<=36'd00000000;
					10'd0847: dataout<=36'd00000000;
					10'd0848: dataout<=36'd00000000;
					10'd0849: dataout<=36'd00000000;
					10'd0850: dataout<=36'd00000000;
					10'd0851: dataout<=36'd00000000;
					10'd0852: dataout<=36'd00000000;
					10'd0853: dataout<=36'd00000000;
					10'd0854: dataout<=36'd00000000;
					10'd0855: dataout<=36'd00000000;
					10'd0856: dataout<=36'd00000000;
					10'd0857: dataout<=36'd00000000;
					10'd0858: dataout<=36'd00000000;
					10'd0859: dataout<=36'd00000000;
					10'd0860: dataout<=36'd00000000;
					10'd0861: dataout<=36'd00000000;
					10'd0862: dataout<=36'd00000000;
					10'd0863: dataout<=36'd00000000;
					10'd0864: dataout<=36'd00000000;
					10'd0865: dataout<=36'd00000000;
					10'd0866: dataout<=36'd00000000;
					10'd0867: dataout<=36'd00000000;
					10'd0868: dataout<=36'd00000000;
					10'd0869: dataout<=36'd00000000;
					10'd0870: dataout<=36'd00000000;
					10'd0871: dataout<=36'd00000000;
					10'd0872: dataout<=36'd00000000;
					10'd0873: dataout<=36'd00000000;
					10'd0874: dataout<=36'd00000000;
					10'd0875: dataout<=36'd00000000;
					10'd0876: dataout<=36'd00000000;
					10'd0877: dataout<=36'd00000000;
					10'd0878: dataout<=36'd00000000;
					10'd0879: dataout<=36'd00000000;
					10'd0880: dataout<=36'd00000000;
					10'd0881: dataout<=36'd00000000;
					10'd0882: dataout<=36'd00000000;
					10'd0883: dataout<=36'd00000000;
					10'd0884: dataout<=36'd00000000;
					10'd0885: dataout<=36'd00000000;
					10'd0886: dataout<=36'd00000000;
					10'd0887: dataout<=36'd00000000;
					10'd0888: dataout<=36'd00000000;
					10'd0889: dataout<=36'd00000000;
					10'd0890: dataout<=36'd00000000;
					10'd0891: dataout<=36'd00000000;
					10'd0892: dataout<=36'd00000000;
					10'd0893: dataout<=36'd00000000;
					10'd0894: dataout<=36'd00000000;
					10'd0895: dataout<=36'd00000000;
					10'd0896: dataout<=36'd00000000;
					10'd0897: dataout<=36'd00000000;
					10'd0898: dataout<=36'd00000000;
					10'd0899: dataout<=36'd00000000;
					10'd0900: dataout<=36'd00000000;
					10'd0901: dataout<=36'd00000000;
					10'd0902: dataout<=36'd00000000;
					10'd0903: dataout<=36'd00000000;
					10'd0904: dataout<=36'd00000000;
					10'd0905: dataout<=36'd00000000;
					10'd0906: dataout<=36'd00000000;
					10'd0907: dataout<=36'd00000000;
					10'd0908: dataout<=36'd00000000;
					10'd0909: dataout<=36'd00000000;
					10'd0910: dataout<=36'd00000000;
					10'd0911: dataout<=36'd00000000;
					10'd0912: dataout<=36'd00000000;
					10'd0913: dataout<=36'd00000000;
					10'd0914: dataout<=36'd00000000;
					10'd0915: dataout<=36'd00000000;
					10'd0916: dataout<=36'd00000000;
					10'd0917: dataout<=36'd00000000;
					10'd0918: dataout<=36'd00000000;
					10'd0919: dataout<=36'd00000000;
					10'd0920: dataout<=36'd00000000;
					10'd0921: dataout<=36'd00000000;
					10'd0922: dataout<=36'd00000000;
					10'd0923: dataout<=36'd00000000;
					10'd0924: dataout<=36'd00000000;
					10'd0925: dataout<=36'd00000000;
					10'd0926: dataout<=36'd00000000;
					10'd0927: dataout<=36'd00000000;
					10'd0928: dataout<=36'd00000000;
					10'd0929: dataout<=36'd00000000;
					10'd0930: dataout<=36'd00000000;
					10'd0931: dataout<=36'd00000000;
					10'd0932: dataout<=36'd00000000;
					10'd0933: dataout<=36'd00000000;
					10'd0934: dataout<=36'd00000000;
					10'd0935: dataout<=36'd00000000;
					10'd0936: dataout<=36'd00000000;
					10'd0937: dataout<=36'd00000000;
					10'd0938: dataout<=36'd00000000;
					10'd0939: dataout<=36'd00000000;
					10'd0940: dataout<=36'd00000000;
					10'd0941: dataout<=36'd00000000;
					10'd0942: dataout<=36'd00000000;
					10'd0943: dataout<=36'd00000000;
					10'd0944: dataout<=36'd00000000;
					10'd0945: dataout<=36'd00000000;
					10'd0946: dataout<=36'd00000000;
					10'd0947: dataout<=36'd00000000;
					10'd0948: dataout<=36'd00000000;
					10'd0949: dataout<=36'd00000000;
					10'd0950: dataout<=36'd00000000;
					10'd0951: dataout<=36'd00000000;
					10'd0952: dataout<=36'd00000000;
					10'd0953: dataout<=36'd00000000;
					10'd0954: dataout<=36'd00000000;
					10'd0955: dataout<=36'd00000000;
					10'd0956: dataout<=36'd00000000;
					10'd0957: dataout<=36'd00000000;
					10'd0958: dataout<=36'd00000000;
					10'd0959: dataout<=36'd00000000;
					10'd0960: dataout<=36'd00000000;
					10'd0961: dataout<=36'd00000000;
					10'd0962: dataout<=36'd00000000;
					10'd0963: dataout<=36'd00000000;
					10'd0964: dataout<=36'd00000000;
					10'd0965: dataout<=36'd00000000;
					10'd0966: dataout<=36'd00000000;
					10'd0967: dataout<=36'd00000000;
					10'd0968: dataout<=36'd00000000;
					10'd0969: dataout<=36'd00000000;
					10'd0970: dataout<=36'd00000000;
					10'd0971: dataout<=36'd00000000;
					10'd0972: dataout<=36'd00000000;
					10'd0973: dataout<=36'd00000000;
					10'd0974: dataout<=36'd00000000;
					10'd0975: dataout<=36'd00000000;
					10'd0976: dataout<=36'd00000000;
					10'd0977: dataout<=36'd00000000;
					10'd0978: dataout<=36'd00000000;
					10'd0979: dataout<=36'd00000000;
					10'd0980: dataout<=36'd00000000;
					10'd0981: dataout<=36'd00000000;
					10'd0982: dataout<=36'd00000000;
					10'd0983: dataout<=36'd00000000;
					10'd0984: dataout<=36'd00000000;
					10'd0985: dataout<=36'd00000000;
					10'd0986: dataout<=36'd00000000;
					10'd0987: dataout<=36'd00000000;
					10'd0988: dataout<=36'd00000000;
					10'd0989: dataout<=36'd00000000;
					10'd0990: dataout<=36'd00000000;
					10'd0991: dataout<=36'd00000000;
					10'd0992: dataout<=36'd00000000;
					10'd0993: dataout<=36'd00000000;
					10'd0994: dataout<=36'd00000000;
					10'd0995: dataout<=36'd00000000;
					10'd0996: dataout<=36'd00000000;
					10'd0997: dataout<=36'd00000000;
					10'd0998: dataout<=36'd00000000;
					10'd0999: dataout<=36'd00000000;
					10'd1000: dataout<=36'd00000000;
					10'd1001: dataout<=36'd00000000;
					10'd1002: dataout<=36'd00000000;
					10'd1003: dataout<=36'd00000000;
					10'd1004: dataout<=36'd00000000;
					10'd1005: dataout<=36'd00000000;
					10'd1006: dataout<=36'd00000000;
					10'd1007: dataout<=36'd00000000;
					10'd1008: dataout<=36'd00000000;
					10'd1009: dataout<=36'd00000000;
					10'd1010: dataout<=36'd00000000;
					10'd1011: dataout<=36'd00000000;
					10'd1012: dataout<=36'd00000000;
					10'd1013: dataout<=36'd00000000;
					10'd1014: dataout<=36'd00000000;
					10'd1015: dataout<=36'd00000000;
					10'd1016: dataout<=36'd00000000;
					10'd1017: dataout<=36'd00000000;
					10'd1018: dataout<=36'd00000000;
					10'd1019: dataout<=36'd00000000;
					10'd1020: dataout<=36'd00000000;
					10'd1021: dataout<=36'd00000000;
					10'd1022: dataout<=36'd00000000;
					10'd1023: dataout<=36'd00000000;
				endcase
			end
		end
	end
endmodule

