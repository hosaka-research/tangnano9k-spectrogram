module nco_rom (clock,ce,oce,reset,addr,dataout);
	input clock,ce,oce,reset;
	input [10:0] addr;
	output [17:0] dataout;
	reg [17:0] dataout;
	always @(posedge clock or posedge reset) begin
		if(reset) begin
			dataout <= 0;
		end else begin
			if (ce & oce) begin
				case (addr)
					11'h0000: dataout<=18'h093fb;
					11'h0001: dataout<=18'h215dc;
					11'h0002: dataout<=18'h264f6;
					11'h0003: dataout<=18'h13143;
					11'h0004: dataout<=18'h08edd;
					11'h0005: dataout<=18'h21457;
					11'h0006: dataout<=18'h2668f;
					11'h0007: dataout<=18'h13367;
					11'h0008: dataout<=18'h089ba;
					11'h0009: dataout<=18'h212e1;
					11'h000a: dataout<=18'h2682b;
					11'h000b: dataout<=18'h13588;
					11'h000c: dataout<=18'h08494;
					11'h000d: dataout<=18'h21178;
					11'h000e: dataout<=18'h269ca;
					11'h000f: dataout<=18'h137a8;
					11'h0010: dataout<=18'h07f6a;
					11'h0011: dataout<=18'h2101d;
					11'h0012: dataout<=18'h26b6b;
					11'h0013: dataout<=18'h139c5;
					11'h0014: dataout<=18'h07a3c;
					11'h0015: dataout<=18'h20ed0;
					11'h0016: dataout<=18'h26d0f;
					11'h0017: dataout<=18'h13be0;
					11'h0018: dataout<=18'h0750b;
					11'h0019: dataout<=18'h20d90;
					11'h001a: dataout<=18'h26eb6;
					11'h001b: dataout<=18'h13df8;
					11'h001c: dataout<=18'h06fd7;
					11'h001d: dataout<=18'h20c5f;
					11'h001e: dataout<=18'h27060;
					11'h001f: dataout<=18'h1400f;
					11'h0020: dataout<=18'h06aa0;
					11'h0021: dataout<=18'h20b3b;
					11'h0022: dataout<=18'h2720d;
					11'h0023: dataout<=18'h14223;
					11'h0024: dataout<=18'h06565;
					11'h0025: dataout<=18'h20a26;
					11'h0026: dataout<=18'h273bc;
					11'h0027: dataout<=18'h14435;
					11'h0028: dataout<=18'h06028;
					11'h0029: dataout<=18'h2091e;
					11'h002a: dataout<=18'h2756e;
					11'h002b: dataout<=18'h14645;
					11'h002c: dataout<=18'h05ae8;
					11'h002d: dataout<=18'h20824;
					11'h002e: dataout<=18'h27723;
					11'h002f: dataout<=18'h14853;
					11'h0030: dataout<=18'h055a6;
					11'h0031: dataout<=18'h20739;
					11'h0032: dataout<=18'h278db;
					11'h0033: dataout<=18'h14a5e;
					11'h0034: dataout<=18'h05061;
					11'h0035: dataout<=18'h2065b;
					11'h0036: dataout<=18'h27a95;
					11'h0037: dataout<=18'h14c67;
					11'h0038: dataout<=18'h04b1a;
					11'h0039: dataout<=18'h2058b;
					11'h003a: dataout<=18'h27c52;
					11'h003b: dataout<=18'h14e6e;
					11'h003c: dataout<=18'h045d1;
					11'h003d: dataout<=18'h204ca;
					11'h003e: dataout<=18'h27e12;
					11'h003f: dataout<=18'h15072;
					11'h0040: dataout<=18'h04086;
					11'h0041: dataout<=18'h20417;
					11'h0042: dataout<=18'h27fd4;
					11'h0043: dataout<=18'h15274;
					11'h0044: dataout<=18'h03b39;
					11'h0045: dataout<=18'h20371;
					11'h0046: dataout<=18'h28199;
					11'h0047: dataout<=18'h15473;
					11'h0048: dataout<=18'h035eb;
					11'h0049: dataout<=18'h202da;
					11'h004a: dataout<=18'h28361;
					11'h004b: dataout<=18'h15671;
					11'h004c: dataout<=18'h0309b;
					11'h004d: dataout<=18'h20252;
					11'h004e: dataout<=18'h2852c;
					11'h004f: dataout<=18'h1586c;
					11'h0050: dataout<=18'h02b4a;
					11'h0051: dataout<=18'h201d7;
					11'h0052: dataout<=18'h286f9;
					11'h0053: dataout<=18'h15a64;
					11'h0054: dataout<=18'h025f7;
					11'h0055: dataout<=18'h2016a;
					11'h0056: dataout<=18'h288c8;
					11'h0057: dataout<=18'h15c5a;
					11'h0058: dataout<=18'h020a4;
					11'h0059: dataout<=18'h2010c;
					11'h005a: dataout<=18'h28a9b;
					11'h005b: dataout<=18'h15e4e;
					11'h005c: dataout<=18'h01b4f;
					11'h005d: dataout<=18'h200bc;
					11'h005e: dataout<=18'h28c70;
					11'h005f: dataout<=18'h1603f;
					11'h0060: dataout<=18'h015fa;
					11'h0061: dataout<=18'h2007a;
					11'h0062: dataout<=18'h28e47;
					11'h0063: dataout<=18'h1622e;
					11'h0064: dataout<=18'h010a4;
					11'h0065: dataout<=18'h20047;
					11'h0066: dataout<=18'h29021;
					11'h0067: dataout<=18'h1641a;
					11'h0068: dataout<=18'h00b4e;
					11'h0069: dataout<=18'h20021;
					11'h006a: dataout<=18'h291fe;
					11'h006b: dataout<=18'h16604;
					11'h006c: dataout<=18'h005f7;
					11'h006d: dataout<=18'h2000a;
					11'h006e: dataout<=18'h293dd;
					11'h006f: dataout<=18'h167eb;
					11'h0070: dataout<=18'h000a0;
					11'h0071: dataout<=18'h20002;
					11'h0072: dataout<=18'h295be;
					11'h0073: dataout<=18'h169d0;
					11'h0074: dataout<=18'h3fb4a;
					11'h0075: dataout<=18'h20007;
					11'h0076: dataout<=18'h297a3;
					11'h0077: dataout<=18'h16bb2;
					11'h0078: dataout<=18'h3f5f4;
					11'h0079: dataout<=18'h2001b;
					11'h007a: dataout<=18'h29989;
					11'h007b: dataout<=18'h16d92;
					11'h007c: dataout<=18'h3f09d;
					11'h007d: dataout<=18'h2003d;
					11'h007e: dataout<=18'h29b73;
					11'h007f: dataout<=18'h16f6f;
					11'h0080: dataout<=18'h3eb47;
					11'h0081: dataout<=18'h2006d;
					11'h0082: dataout<=18'h29d5e;
					11'h0083: dataout<=18'h1714a;
					11'h0084: dataout<=18'h3e5f2;
					11'h0085: dataout<=18'h200ab;
					11'h0086: dataout<=18'h29f4c;
					11'h0087: dataout<=18'h17322;
					11'h0088: dataout<=18'h3e09d;
					11'h0089: dataout<=18'h200f8;
					11'h008a: dataout<=18'h2a13d;
					11'h008b: dataout<=18'h174f7;
					11'h008c: dataout<=18'h3db4a;
					11'h008d: dataout<=18'h20153;
					11'h008e: dataout<=18'h2a330;
					11'h008f: dataout<=18'h176ca;
					11'h0090: dataout<=18'h3d5f7;
					11'h0091: dataout<=18'h201bc;
					11'h0092: dataout<=18'h2a526;
					11'h0093: dataout<=18'h1789a;
					11'h0094: dataout<=18'h3d0a5;
					11'h0095: dataout<=18'h20233;
					11'h0096: dataout<=18'h2a71e;
					11'h0097: dataout<=18'h17a68;
					11'h0098: dataout<=18'h3cb55;
					11'h0099: dataout<=18'h202b9;
					11'h009a: dataout<=18'h2a918;
					11'h009b: dataout<=18'h17c33;
					11'h009c: dataout<=18'h3c606;
					11'h009d: dataout<=18'h2034d;
					11'h009e: dataout<=18'h2ab15;
					11'h009f: dataout<=18'h17dfc;
					11'h00a0: dataout<=18'h3c0b9;
					11'h00a1: dataout<=18'h203ee;
					11'h00a2: dataout<=18'h2ad14;
					11'h00a3: dataout<=18'h17fc1;
					11'h00a4: dataout<=18'h3bb6d;
					11'h00a5: dataout<=18'h2049e;
					11'h00a6: dataout<=18'h2af15;
					11'h00a7: dataout<=18'h18184;
					11'h00a8: dataout<=18'h3b624;
					11'h00a9: dataout<=18'h2055d;
					11'h00aa: dataout<=18'h2b119;
					11'h00ab: dataout<=18'h18345;
					11'h00ac: dataout<=18'h3b0dc;
					11'h00ad: dataout<=18'h20629;
					11'h00ae: dataout<=18'h2b31f;
					11'h00af: dataout<=18'h18502;
					11'h00b0: dataout<=18'h3ab97;
					11'h00b1: dataout<=18'h20703;
					11'h00b2: dataout<=18'h2b527;
					11'h00b3: dataout<=18'h186bd;
					11'h00b4: dataout<=18'h3a654;
					11'h00b5: dataout<=18'h207eb;
					11'h00b6: dataout<=18'h2b732;
					11'h00b7: dataout<=18'h18876;
					11'h00b8: dataout<=18'h3a114;
					11'h00b9: dataout<=18'h208e2;
					11'h00ba: dataout<=18'h2b93f;
					11'h00bb: dataout<=18'h18a2b;
					11'h00bc: dataout<=18'h39bd6;
					11'h00bd: dataout<=18'h209e6;
					11'h00be: dataout<=18'h2bb4e;
					11'h00bf: dataout<=18'h18bde;
					11'h00c0: dataout<=18'h3969b;
					11'h00c1: dataout<=18'h20af9;
					11'h00c2: dataout<=18'h2bd60;
					11'h00c3: dataout<=18'h18d8e;
					11'h00c4: dataout<=18'h39163;
					11'h00c5: dataout<=18'h20c19;
					11'h00c6: dataout<=18'h2bf74;
					11'h00c7: dataout<=18'h18f3b;
					11'h00c8: dataout<=18'h38c2e;
					11'h00c9: dataout<=18'h20d47;
					11'h00ca: dataout<=18'h2c18a;
					11'h00cb: dataout<=18'h190e6;
					11'h00cc: dataout<=18'h386fc;
					11'h00cd: dataout<=18'h20e83;
					11'h00ce: dataout<=18'h2c3a2;
					11'h00cf: dataout<=18'h1928d;
					11'h00d0: dataout<=18'h381ce;
					11'h00d1: dataout<=18'h20fcd;
					11'h00d2: dataout<=18'h2c5bc;
					11'h00d3: dataout<=18'h19432;
					11'h00d4: dataout<=18'h37ca3;
					11'h00d5: dataout<=18'h21125;
					11'h00d6: dataout<=18'h2c7d9;
					11'h00d7: dataout<=18'h195d4;
					11'h00d8: dataout<=18'h3777c;
					11'h00d9: dataout<=18'h2128b;
					11'h00da: dataout<=18'h2c9f8;
					11'h00db: dataout<=18'h19774;
					11'h00dc: dataout<=18'h37258;
					11'h00dd: dataout<=18'h213fe;
					11'h00de: dataout<=18'h2cc19;
					11'h00df: dataout<=18'h19910;
					11'h00e0: dataout<=18'h36d39;
					11'h00e1: dataout<=18'h2157f;
					11'h00e2: dataout<=18'h2ce3c;
					11'h00e3: dataout<=18'h19aaa;
					11'h00e4: dataout<=18'h3681d;
					11'h00e5: dataout<=18'h2170e;
					11'h00e6: dataout<=18'h2d061;
					11'h00e7: dataout<=18'h19c40;
					11'h00e8: dataout<=18'h36306;
					11'h00e9: dataout<=18'h218aa;
					11'h00ea: dataout<=18'h2d288;
					11'h00eb: dataout<=18'h19dd4;
					11'h00ec: dataout<=18'h35df3;
					11'h00ed: dataout<=18'h21a54;
					11'h00ee: dataout<=18'h2d4b2;
					11'h00ef: dataout<=18'h19f65;
					11'h00f0: dataout<=18'h358e5;
					11'h00f1: dataout<=18'h21c0b;
					11'h00f2: dataout<=18'h2d6dd;
					11'h00f3: dataout<=18'h1a0f3;
					11'h00f4: dataout<=18'h353dc;
					11'h00f5: dataout<=18'h21dd0;
					11'h00f6: dataout<=18'h2d90b;
					11'h00f7: dataout<=18'h1a27e;
					11'h00f8: dataout<=18'h34ed7;
					11'h00f9: dataout<=18'h21fa2;
					11'h00fa: dataout<=18'h2db3a;
					11'h00fb: dataout<=18'h1a407;
					11'h00fc: dataout<=18'h349d7;
					11'h00fd: dataout<=18'h22182;
					11'h00fe: dataout<=18'h2dd6c;
					11'h00ff: dataout<=18'h1a58c;
					11'h0100: dataout<=18'h344dc;
					11'h0101: dataout<=18'h2236f;
					11'h0102: dataout<=18'h2dfa0;
					11'h0103: dataout<=18'h1a70e;
					11'h0104: dataout<=18'h33fe6;
					11'h0105: dataout<=18'h22569;
					11'h0106: dataout<=18'h2e1d5;
					11'h0107: dataout<=18'h1a88e;
					11'h0108: dataout<=18'h33af6;
					11'h0109: dataout<=18'h22771;
					11'h010a: dataout<=18'h2e40d;
					11'h010b: dataout<=18'h1aa0a;
					11'h010c: dataout<=18'h3360b;
					11'h010d: dataout<=18'h22985;
					11'h010e: dataout<=18'h2e647;
					11'h010f: dataout<=18'h1ab84;
					11'h0110: dataout<=18'h33126;
					11'h0111: dataout<=18'h22ba7;
					11'h0112: dataout<=18'h2e882;
					11'h0113: dataout<=18'h1acfa;
					11'h0114: dataout<=18'h32c47;
					11'h0115: dataout<=18'h22dd6;
					11'h0116: dataout<=18'h2eac0;
					11'h0117: dataout<=18'h1ae6e;
					11'h0118: dataout<=18'h3276d;
					11'h0119: dataout<=18'h23011;
					11'h011a: dataout<=18'h2ed00;
					11'h011b: dataout<=18'h1afdf;
					11'h011c: dataout<=18'h3229a;
					11'h011d: dataout<=18'h2325a;
					11'h011e: dataout<=18'h2ef41;
					11'h011f: dataout<=18'h1b14c;
					11'h0120: dataout<=18'h31dcc;
					11'h0121: dataout<=18'h234af;
					11'h0122: dataout<=18'h2f184;
					11'h0123: dataout<=18'h1b2b7;
					11'h0124: dataout<=18'h31905;
					11'h0125: dataout<=18'h23712;
					11'h0126: dataout<=18'h2f3c9;
					11'h0127: dataout<=18'h1b41e;
					11'h0128: dataout<=18'h31445;
					11'h0129: dataout<=18'h23981;
					11'h012a: dataout<=18'h2f611;
					11'h012b: dataout<=18'h1b583;
					11'h012c: dataout<=18'h30f8b;
					11'h012d: dataout<=18'h23bfc;
					11'h012e: dataout<=18'h2f859;
					11'h012f: dataout<=18'h1b6e4;
					11'h0130: dataout<=18'h30ad7;
					11'h0131: dataout<=18'h23e84;
					11'h0132: dataout<=18'h2faa4;
					11'h0133: dataout<=18'h1b843;
					11'h0134: dataout<=18'h3062b;
					11'h0135: dataout<=18'h24119;
					11'h0136: dataout<=18'h2fcf1;
					11'h0137: dataout<=18'h1b99e;
					11'h0138: dataout<=18'h30185;
					11'h0139: dataout<=18'h243ba;
					11'h013a: dataout<=18'h2ff3f;
					11'h013b: dataout<=18'h1baf6;
					11'h013c: dataout<=18'h2fce7;
					11'h013d: dataout<=18'h24668;
					11'h013e: dataout<=18'h3018f;
					11'h013f: dataout<=18'h1bc4b;
					11'h0140: dataout<=18'h2f850;
					11'h0141: dataout<=18'h24922;
					11'h0142: dataout<=18'h303e1;
					11'h0143: dataout<=18'h1bd9d;
					11'h0144: dataout<=18'h2f3c0;
					11'h0145: dataout<=18'h24be8;
					11'h0146: dataout<=18'h30635;
					11'h0147: dataout<=18'h1beec;
					11'h0148: dataout<=18'h2ef37;
					11'h0149: dataout<=18'h24eba;
					11'h014a: dataout<=18'h3088a;
					11'h014b: dataout<=18'h1c038;
					11'h014c: dataout<=18'h2eab6;
					11'h014d: dataout<=18'h25198;
					11'h014e: dataout<=18'h30ae1;
					11'h014f: dataout<=18'h1c181;
					11'h0150: dataout<=18'h2e63d;
					11'h0151: dataout<=18'h25482;
					11'h0152: dataout<=18'h30d3a;
					11'h0153: dataout<=18'h1c2c7;
					11'h0154: dataout<=18'h2e1cc;
					11'h0155: dataout<=18'h25779;
					11'h0156: dataout<=18'h30f95;
					11'h0157: dataout<=18'h1c409;
					11'h0158: dataout<=18'h2dd63;
					11'h0159: dataout<=18'h25a7b;
					11'h015a: dataout<=18'h311f1;
					11'h015b: dataout<=18'h1c548;
					11'h015c: dataout<=18'h2d901;
					11'h015d: dataout<=18'h25d88;
					11'h015e: dataout<=18'h3144f;
					11'h015f: dataout<=18'h1c685;
					11'h0160: dataout<=18'h2d4a8;
					11'h0161: dataout<=18'h260a2;
					11'h0162: dataout<=18'h316ae;
					11'h0163: dataout<=18'h1c7be;
					11'h0164: dataout<=18'h2d058;
					11'h0165: dataout<=18'h263c6;
					11'h0166: dataout<=18'h31910;
					11'h0167: dataout<=18'h1c8f4;
					11'h0168: dataout<=18'h2cc0f;
					11'h0169: dataout<=18'h266f7;
					11'h016a: dataout<=18'h31b72;
					11'h016b: dataout<=18'h1ca26;
					11'h016c: dataout<=18'h2c7d0;
					11'h016d: dataout<=18'h26a33;
					11'h016e: dataout<=18'h31dd7;
					11'h016f: dataout<=18'h1cb56;
					11'h0170: dataout<=18'h2c399;
					11'h0171: dataout<=18'h26d7a;
					11'h0172: dataout<=18'h3203d;
					11'h0173: dataout<=18'h1cc82;
					11'h0174: dataout<=18'h2bf6b;
					11'h0175: dataout<=18'h270cc;
					11'h0176: dataout<=18'h322a4;
					11'h0177: dataout<=18'h1cdab;
					11'h0178: dataout<=18'h2bb45;
					11'h0179: dataout<=18'h27429;
					11'h017a: dataout<=18'h3250d;
					11'h017b: dataout<=18'h1ced1;
					11'h017c: dataout<=18'h2b729;
					11'h017d: dataout<=18'h27792;
					11'h017e: dataout<=18'h32778;
					11'h017f: dataout<=18'h1cff4;
					11'h0180: dataout<=18'h2b316;
					11'h0181: dataout<=18'h27b05;
					11'h0182: dataout<=18'h329e4;
					11'h0183: dataout<=18'h1d113;
					11'h0184: dataout<=18'h2af0c;
					11'h0185: dataout<=18'h27e83;
					11'h0186: dataout<=18'h32c51;
					11'h0187: dataout<=18'h1d22f;
					11'h0188: dataout<=18'h2ab0c;
					11'h0189: dataout<=18'h2820c;
					11'h018a: dataout<=18'h32ec0;
					11'h018b: dataout<=18'h1d348;
					11'h018c: dataout<=18'h2a715;
					11'h018d: dataout<=18'h285a0;
					11'h018e: dataout<=18'h33131;
					11'h018f: dataout<=18'h1d45e;
					11'h0190: dataout<=18'h2a328;
					11'h0191: dataout<=18'h2893e;
					11'h0192: dataout<=18'h333a3;
					11'h0193: dataout<=18'h1d570;
					11'h0194: dataout<=18'h29f44;
					11'h0195: dataout<=18'h28ce6;
					11'h0196: dataout<=18'h33616;
					11'h0197: dataout<=18'h1d67f;
					11'h0198: dataout<=18'h29b6a;
					11'h0199: dataout<=18'h29099;
					11'h019a: dataout<=18'h3388b;
					11'h019b: dataout<=18'h1d78b;
					11'h019c: dataout<=18'h2979b;
					11'h019d: dataout<=18'h29456;
					11'h019e: dataout<=18'h33b01;
					11'h019f: dataout<=18'h1d894;
					11'h01a0: dataout<=18'h293d5;
					11'h01a1: dataout<=18'h2981d;
					11'h01a2: dataout<=18'h33d78;
					11'h01a3: dataout<=18'h1d999;
					11'h01a4: dataout<=18'h29019;
					11'h01a5: dataout<=18'h29bee;
					11'h01a6: dataout<=18'h33ff1;
					11'h01a7: dataout<=18'h1da9b;
					11'h01a8: dataout<=18'h28c68;
					11'h01a9: dataout<=18'h29fc9;
					11'h01aa: dataout<=18'h3426b;
					11'h01ab: dataout<=18'h1db9a;
					11'h01ac: dataout<=18'h288c1;
					11'h01ad: dataout<=18'h2a3ae;
					11'h01ae: dataout<=18'h344e7;
					11'h01af: dataout<=18'h1dc95;
					11'h01b0: dataout<=18'h28524;
					11'h01b1: dataout<=18'h2a79d;
					11'h01b2: dataout<=18'h34763;
					11'h01b3: dataout<=18'h1dd8d;
					11'h01b4: dataout<=18'h28192;
					11'h01b5: dataout<=18'h2ab95;
					11'h01b6: dataout<=18'h349e2;
					11'h01b7: dataout<=18'h1de82;
					11'h01b8: dataout<=18'h27e0a;
					11'h01b9: dataout<=18'h2af97;
					11'h01ba: dataout<=18'h34c61;
					11'h01bb: dataout<=18'h1df74;
					11'h01bc: dataout<=18'h27a8e;
					11'h01bd: dataout<=18'h2b3a2;
					11'h01be: dataout<=18'h34ee1;
					11'h01bf: dataout<=18'h1e062;
					11'h01c0: dataout<=18'h2771c;
					11'h01c1: dataout<=18'h2b7b6;
					11'h01c2: dataout<=18'h35163;
					11'h01c3: dataout<=18'h1e14c;
					11'h01c4: dataout<=18'h273b5;
					11'h01c5: dataout<=18'h2bbd4;
					11'h01c6: dataout<=18'h353e6;
					11'h01c7: dataout<=18'h1e234;
					11'h01c8: dataout<=18'h27059;
					11'h01c9: dataout<=18'h2bffa;
					11'h01ca: dataout<=18'h3566b;
					11'h01cb: dataout<=18'h1e318;
					11'h01cc: dataout<=18'h26d08;
					11'h01cd: dataout<=18'h2c429;
					11'h01ce: dataout<=18'h358f0;
					11'h01cf: dataout<=18'h1e3f8;
					11'h01d0: dataout<=18'h269c3;
					11'h01d1: dataout<=18'h2c861;
					11'h01d2: dataout<=18'h35b77;
					11'h01d3: dataout<=18'h1e4d6;
					11'h01d4: dataout<=18'h26688;
					11'h01d5: dataout<=18'h2cca2;
					11'h01d6: dataout<=18'h35dfe;
					11'h01d7: dataout<=18'h1e5b0;
					11'h01d8: dataout<=18'h2635a;
					11'h01d9: dataout<=18'h2d0ec;
					11'h01da: dataout<=18'h36087;
					11'h01db: dataout<=18'h1e686;
					11'h01dc: dataout<=18'h26036;
					11'h01dd: dataout<=18'h2d53e;
					11'h01de: dataout<=18'h36311;
					11'h01df: dataout<=18'h1e759;
					11'h01e0: dataout<=18'h25d1e;
					11'h01e1: dataout<=18'h2d998;
					11'h01e2: dataout<=18'h3659c;
					11'h01e3: dataout<=18'h1e829;
					11'h01e4: dataout<=18'h25a12;
					11'h01e5: dataout<=18'h2ddfa;
					11'h01e6: dataout<=18'h36828;
					11'h01e7: dataout<=18'h1e8f6;
					11'h01e8: dataout<=18'h25712;
					11'h01e9: dataout<=18'h2e264;
					11'h01ea: dataout<=18'h36ab6;
					11'h01eb: dataout<=18'h1e9bf;
					11'h01ec: dataout<=18'h2541d;
					11'h01ed: dataout<=18'h2e6d7;
					11'h01ee: dataout<=18'h36d44;
					11'h01ef: dataout<=18'h1ea84;
					11'h01f0: dataout<=18'h25135;
					11'h01f1: dataout<=18'h2eb51;
					11'h01f2: dataout<=18'h36fd3;
					11'h01f3: dataout<=18'h1eb46;
					11'h01f4: dataout<=18'h24e58;
					11'h01f5: dataout<=18'h2efd3;
					11'h01f6: dataout<=18'h37263;
					11'h01f7: dataout<=18'h1ec05;
					11'h01f8: dataout<=18'h24b88;
					11'h01f9: dataout<=18'h2f45c;
					11'h01fa: dataout<=18'h374f5;
					11'h01fb: dataout<=18'h1ecc0;
					11'h01fc: dataout<=18'h248c3;
					11'h01fd: dataout<=18'h2f8ed;
					11'h01fe: dataout<=18'h37787;
					11'h01ff: dataout<=18'h1ed78;
					11'h0200: dataout<=18'h2460b;
					11'h0201: dataout<=18'h2fd85;
					11'h0202: dataout<=18'h37a1a;
					11'h0203: dataout<=18'h1ee2d;
					11'h0204: dataout<=18'h2435f;
					11'h0205: dataout<=18'h30225;
					11'h0206: dataout<=18'h37cae;
					11'h0207: dataout<=18'h1eede;
					11'h0208: dataout<=18'h240c0;
					11'h0209: dataout<=18'h306cb;
					11'h020a: dataout<=18'h37f43;
					11'h020b: dataout<=18'h1ef8b;
					11'h020c: dataout<=18'h23e2d;
					11'h020d: dataout<=18'h30b79;
					11'h020e: dataout<=18'h381d9;
					11'h020f: dataout<=18'h1f035;
					11'h0210: dataout<=18'h23ba6;
					11'h0211: dataout<=18'h3102d;
					11'h0212: dataout<=18'h38470;
					11'h0213: dataout<=18'h1f0dc;
					11'h0214: dataout<=18'h2392c;
					11'h0215: dataout<=18'h314e8;
					11'h0216: dataout<=18'h38707;
					11'h0217: dataout<=18'h1f17f;
					11'h0218: dataout<=18'h236bf;
					11'h0219: dataout<=18'h319a9;
					11'h021a: dataout<=18'h389a0;
					11'h021b: dataout<=18'h1f21f;
					11'h021c: dataout<=18'h2345e;
					11'h021d: dataout<=18'h31e71;
					11'h021e: dataout<=18'h38c39;
					11'h021f: dataout<=18'h1f2bb;
					11'h0220: dataout<=18'h2320b;
					11'h0221: dataout<=18'h3233f;
					11'h0222: dataout<=18'h38ed3;
					11'h0223: dataout<=18'h1f354;
					11'h0224: dataout<=18'h22fc4;
					11'h0225: dataout<=18'h32814;
					11'h0226: dataout<=18'h3916e;
					11'h0227: dataout<=18'h1f3e9;
					11'h0228: dataout<=18'h22d8a;
					11'h0229: dataout<=18'h32cee;
					11'h022a: dataout<=18'h3940a;
					11'h022b: dataout<=18'h1f47b;
					11'h022c: dataout<=18'h22b5d;
					11'h022d: dataout<=18'h331ce;
					11'h022e: dataout<=18'h396a6;
					11'h022f: dataout<=18'h1f50a;
					11'h0230: dataout<=18'h2293d;
					11'h0231: dataout<=18'h336b4;
					11'h0232: dataout<=18'h39943;
					11'h0233: dataout<=18'h1f595;
					11'h0234: dataout<=18'h2272a;
					11'h0235: dataout<=18'h33ba0;
					11'h0236: dataout<=18'h39be1;
					11'h0237: dataout<=18'h1f61c;
					11'h0238: dataout<=18'h22524;
					11'h0239: dataout<=18'h34091;
					11'h023a: dataout<=18'h39e80;
					11'h023b: dataout<=18'h1f6a0;
					11'h023c: dataout<=18'h2232c;
					11'h023d: dataout<=18'h34587;
					11'h023e: dataout<=18'h3a11f;
					11'h023f: dataout<=18'h1f720;
					11'h0240: dataout<=18'h22141;
					11'h0241: dataout<=18'h34a83;
					11'h0242: dataout<=18'h3a3bf;
					11'h0243: dataout<=18'h1f79d;
					11'h0244: dataout<=18'h21f63;
					11'h0245: dataout<=18'h34f83;
					11'h0246: dataout<=18'h3a660;
					11'h0247: dataout<=18'h1f817;
					11'h0248: dataout<=18'h21d92;
					11'h0249: dataout<=18'h35489;
					11'h024a: dataout<=18'h3a901;
					11'h024b: dataout<=18'h1f88c;
					11'h024c: dataout<=18'h21bcf;
					11'h024d: dataout<=18'h35993;
					11'h024e: dataout<=18'h3aba2;
					11'h024f: dataout<=18'h1f8ff;
					11'h0250: dataout<=18'h21a1a;
					11'h0251: dataout<=18'h35ea2;
					11'h0252: dataout<=18'h3ae45;
					11'h0253: dataout<=18'h1f96e;
					11'h0254: dataout<=18'h21872;
					11'h0255: dataout<=18'h363b5;
					11'h0256: dataout<=18'h3b0e8;
					11'h0257: dataout<=18'h1f9d9;
					11'h0258: dataout<=18'h216d7;
					11'h0259: dataout<=18'h368cd;
					11'h025a: dataout<=18'h3b38b;
					11'h025b: dataout<=18'h1fa41;
					11'h025c: dataout<=18'h2154b;
					11'h025d: dataout<=18'h36de9;
					11'h025e: dataout<=18'h3b62f;
					11'h025f: dataout<=18'h1faa5;
					11'h0260: dataout<=18'h213cb;
					11'h0261: dataout<=18'h37309;
					11'h0262: dataout<=18'h3b8d4;
					11'h0263: dataout<=18'h1fb06;
					11'h0264: dataout<=18'h2125a;
					11'h0265: dataout<=18'h3782d;
					11'h0266: dataout<=18'h3bb79;
					11'h0267: dataout<=18'h1fb63;
					11'h0268: dataout<=18'h210f6;
					11'h0269: dataout<=18'h37d55;
					11'h026a: dataout<=18'h3be1e;
					11'h026b: dataout<=18'h1fbbd;
					11'h026c: dataout<=18'h20fa0;
					11'h026d: dataout<=18'h38280;
					11'h026e: dataout<=18'h3c0c4;
					11'h026f: dataout<=18'h1fc13;
					11'h0270: dataout<=18'h20e58;
					11'h0271: dataout<=18'h387af;
					11'h0272: dataout<=18'h3c36b;
					11'h0273: dataout<=18'h1fc66;
					11'h0274: dataout<=18'h20d1e;
					11'h0275: dataout<=18'h38ce1;
					11'h0276: dataout<=18'h3c611;
					11'h0277: dataout<=18'h1fcb5;
					11'h0278: dataout<=18'h20bf1;
					11'h0279: dataout<=18'h39216;
					11'h027a: dataout<=18'h3c8b9;
					11'h027b: dataout<=18'h1fd00;
					11'h027c: dataout<=18'h20ad3;
					11'h027d: dataout<=18'h3974f;
					11'h027e: dataout<=18'h3cb60;
					11'h027f: dataout<=18'h1fd48;
					11'h0280: dataout<=18'h209c2;
					11'h0281: dataout<=18'h39c8a;
					11'h0282: dataout<=18'h3ce08;
					11'h0283: dataout<=18'h1fd8d;
					11'h0284: dataout<=18'h208c0;
					11'h0285: dataout<=18'h3a1c8;
					11'h0286: dataout<=18'h3d0b1;
					11'h0287: dataout<=18'h1fdce;
					11'h0288: dataout<=18'h207cb;
					11'h0289: dataout<=18'h3a709;
					11'h028a: dataout<=18'h3d359;
					11'h028b: dataout<=18'h1fe0b;
					11'h028c: dataout<=18'h206e5;
					11'h028d: dataout<=18'h3ac4c;
					11'h028e: dataout<=18'h3d602;
					11'h028f: dataout<=18'h1fe45;
					11'h0290: dataout<=18'h2060d;
					11'h0291: dataout<=18'h3b192;
					11'h0292: dataout<=18'h3d8ab;
					11'h0293: dataout<=18'h1fe7b;
					11'h0294: dataout<=18'h20542;
					11'h0295: dataout<=18'h3b6da;
					11'h0296: dataout<=18'h3db55;
					11'h0297: dataout<=18'h1feae;
					11'h0298: dataout<=18'h20486;
					11'h0299: dataout<=18'h3bc24;
					11'h029a: dataout<=18'h3ddff;
					11'h029b: dataout<=18'h1fedd;
					11'h029c: dataout<=18'h203d8;
					11'h029d: dataout<=18'h3c16f;
					11'h029e: dataout<=18'h3e0a9;
					11'h029f: dataout<=18'h1ff09;
					11'h02a0: dataout<=18'h20338;
					11'h02a1: dataout<=18'h3c6bd;
					11'h02a2: dataout<=18'h3e353;
					11'h02a3: dataout<=18'h1ff31;
					11'h02a4: dataout<=18'h202a6;
					11'h02a5: dataout<=18'h3cc0c;
					11'h02a6: dataout<=18'h3e5fe;
					11'h02a7: dataout<=18'h1ff55;
					11'h02a8: dataout<=18'h20223;
					11'h02a9: dataout<=18'h3d15c;
					11'h02aa: dataout<=18'h3e8a8;
					11'h02ab: dataout<=18'h1ff76;
					11'h02ac: dataout<=18'h201ad;
					11'h02ad: dataout<=18'h3d6ae;
					11'h02ae: dataout<=18'h3eb53;
					11'h02af: dataout<=18'h1ff94;
					11'h02b0: dataout<=18'h20146;
					11'h02b1: dataout<=18'h3dc01;
					11'h02b2: dataout<=18'h3edfe;
					11'h02b3: dataout<=18'h1ffad;
					11'h02b4: dataout<=18'h200ed;
					11'h02b5: dataout<=18'h3e155;
					11'h02b6: dataout<=18'h3f0a9;
					11'h02b7: dataout<=18'h1ffc4;
					11'h02b8: dataout<=18'h200a2;
					11'h02b9: dataout<=18'h3e6aa;
					11'h02ba: dataout<=18'h3f354;
					11'h02bb: dataout<=18'h1ffd6;
					11'h02bc: dataout<=18'h20066;
					11'h02bd: dataout<=18'h3ebff;
					11'h02be: dataout<=18'h3f5ff;
					11'h02bf: dataout<=18'h1ffe5;
					11'h02c0: dataout<=18'h20037;
					11'h02c1: dataout<=18'h3f155;
					11'h02c2: dataout<=18'h3f8ab;
					11'h02c3: dataout<=18'h1fff1;
					11'h02c4: dataout<=18'h20017;
					11'h02c5: dataout<=18'h3f6ac;
					11'h02c6: dataout<=18'h3fb56;
					11'h02c7: dataout<=18'h1fff9;
					11'h02c8: dataout<=18'h20005;
					11'h02c9: dataout<=18'h3fc02;
					11'h02ca: dataout<=18'h3fe01;
					11'h02cb: dataout<=18'h1fffe;
					11'h02cc: dataout<=18'h20002;
					11'h02cd: dataout<=18'h00158;
					11'h02ce: dataout<=18'h000ac;
					11'h02cf: dataout<=18'h1fffe;
					11'h02d0: dataout<=18'h2000d;
					11'h02d1: dataout<=18'h006af;
					11'h02d2: dataout<=18'h00357;
					11'h02d3: dataout<=18'h1fffc;
					11'h02d4: dataout<=18'h20026;
					11'h02d5: dataout<=18'h00c05;
					11'h02d6: dataout<=18'h00603;
					11'h02d7: dataout<=18'h1fff5;
					11'h02d8: dataout<=18'h2004d;
					11'h02d9: dataout<=18'h0115c;
					11'h02da: dataout<=18'h008ae;
					11'h02db: dataout<=18'h1ffec;
					11'h02dc: dataout<=18'h20082;
					11'h02dd: dataout<=18'h016b1;
					11'h02de: dataout<=18'h00b59;
					11'h02df: dataout<=18'h1ffde;
					11'h02e0: dataout<=18'h200c6;
					11'h02e1: dataout<=18'h01c07;
					11'h02e2: dataout<=18'h00e04;
					11'h02e3: dataout<=18'h1ffcd;
					11'h02e4: dataout<=18'h20118;
					11'h02e5: dataout<=18'h0215b;
					11'h02e6: dataout<=18'h010b0;
					11'h02e7: dataout<=18'h1ffb9;
					11'h02e8: dataout<=18'h20178;
					11'h02e9: dataout<=18'h026ae;
					11'h02ea: dataout<=18'h0135b;
					11'h02eb: dataout<=18'h1ffa1;
					11'h02ec: dataout<=18'h201e7;
					11'h02ed: dataout<=18'h02c01;
					11'h02ee: dataout<=18'h01605;
					11'h02ef: dataout<=18'h1ff85;
					11'h02f0: dataout<=18'h20263;
					11'h02f1: dataout<=18'h03152;
					11'h02f2: dataout<=18'h018b0;
					11'h02f3: dataout<=18'h1ff66;
					11'h02f4: dataout<=18'h202ee;
					11'h02f5: dataout<=18'h036a2;
					11'h02f6: dataout<=18'h01b5b;
					11'h02f7: dataout<=18'h1ff43;
					11'h02f8: dataout<=18'h20387;
					11'h02f9: dataout<=18'h03bf0;
					11'h02fa: dataout<=18'h01e05;
					11'h02fb: dataout<=18'h1ff1d;
					11'h02fc: dataout<=18'h2042e;
					11'h02fd: dataout<=18'h0413d;
					11'h02fe: dataout<=18'h020af;
					11'h02ff: dataout<=18'h1fef3;
					11'h0300: dataout<=18'h204e3;
					11'h0301: dataout<=18'h04687;
					11'h0302: dataout<=18'h02359;
					11'h0303: dataout<=18'h1fec6;
					11'h0304: dataout<=18'h205a6;
					11'h0305: dataout<=18'h04bd0;
					11'h0306: dataout<=18'h02603;
					11'h0307: dataout<=18'h1fe95;
					11'h0308: dataout<=18'h20678;
					11'h0309: dataout<=18'h05117;
					11'h030a: dataout<=18'h028ac;
					11'h030b: dataout<=18'h1fe60;
					11'h030c: dataout<=18'h20757;
					11'h030d: dataout<=18'h0565b;
					11'h030e: dataout<=18'h02b55;
					11'h030f: dataout<=18'h1fe28;
					11'h0310: dataout<=18'h20845;
					11'h0311: dataout<=18'h05b9d;
					11'h0312: dataout<=18'h02dfe;
					11'h0313: dataout<=18'h1fded;
					11'h0314: dataout<=18'h20941;
					11'h0315: dataout<=18'h060dd;
					11'h0316: dataout<=18'h030a6;
					11'h0317: dataout<=18'h1fdad;
					11'h0318: dataout<=18'h20a4a;
					11'h0319: dataout<=18'h06619;
					11'h031a: dataout<=18'h0334f;
					11'h031b: dataout<=18'h1fd6b;
					11'h031c: dataout<=18'h20b62;
					11'h031d: dataout<=18'h06b53;
					11'h031e: dataout<=18'h035f6;
					11'h031f: dataout<=18'h1fd24;
					11'h0320: dataout<=18'h20c87;
					11'h0321: dataout<=18'h0708a;
					11'h0322: dataout<=18'h0389e;
					11'h0323: dataout<=18'h1fcdb;
					11'h0324: dataout<=18'h20dbb;
					11'h0325: dataout<=18'h075be;
					11'h0326: dataout<=18'h03b45;
					11'h0327: dataout<=18'h1fc8d;
					11'h0328: dataout<=18'h20efc;
					11'h0329: dataout<=18'h07aef;
					11'h032a: dataout<=18'h03deb;
					11'h032b: dataout<=18'h1fc3c;
					11'h032c: dataout<=18'h2104b;
					11'h032d: dataout<=18'h0801c;
					11'h032e: dataout<=18'h04092;
					11'h032f: dataout<=18'h1fbe8;
					11'h0330: dataout<=18'h211a8;
					11'h0331: dataout<=18'h08545;
					11'h0332: dataout<=18'h04337;
					11'h0333: dataout<=18'h1fb90;
					11'h0334: dataout<=18'h21312;
					11'h0335: dataout<=18'h08a6b;
					11'h0336: dataout<=18'h045dd;
					11'h0337: dataout<=18'h1fb35;
					11'h0338: dataout<=18'h2148b;
					11'h0339: dataout<=18'h08f8d;
					11'h033a: dataout<=18'h04881;
					11'h033b: dataout<=18'h1fad6;
					11'h033c: dataout<=18'h21611;
					11'h033d: dataout<=18'h094ab;
					11'h033e: dataout<=18'h04b26;
					11'h033f: dataout<=18'h1fa73;
					11'h0340: dataout<=18'h217a5;
					11'h0341: dataout<=18'h099c5;
					11'h0342: dataout<=18'h04dc9;
					11'h0343: dataout<=18'h1fa0d;
					11'h0344: dataout<=18'h21946;
					11'h0345: dataout<=18'h09eda;
					11'h0346: dataout<=18'h0506d;
					11'h0347: dataout<=18'h1f9a3;
					11'h0348: dataout<=18'h21af5;
					11'h0349: dataout<=18'h0a3ec;
					11'h034a: dataout<=18'h0530f;
					11'h034b: dataout<=18'h1f936;
					11'h034c: dataout<=18'h21cb1;
					11'h034d: dataout<=18'h0a8f8;
					11'h034e: dataout<=18'h055b1;
					11'h034f: dataout<=18'h1f8c6;
					11'h0350: dataout<=18'h21e7b;
					11'h0351: dataout<=18'h0ae00;
					11'h0352: dataout<=18'h05853;
					11'h0353: dataout<=18'h1f851;
					11'h0354: dataout<=18'h22052;
					11'h0355: dataout<=18'h0b303;
					11'h0356: dataout<=18'h05af4;
					11'h0357: dataout<=18'h1f7da;
					11'h0358: dataout<=18'h22237;
					11'h0359: dataout<=18'h0b801;
					11'h035a: dataout<=18'h05d94;
					11'h035b: dataout<=18'h1f75f;
					11'h035c: dataout<=18'h22429;
					11'h035d: dataout<=18'h0bcfa;
					11'h035e: dataout<=18'h06033;
					11'h035f: dataout<=18'h1f6e0;
					11'h0360: dataout<=18'h22628;
					11'h0361: dataout<=18'h0c1ee;
					11'h0362: dataout<=18'h062d2;
					11'h0363: dataout<=18'h1f65e;
					11'h0364: dataout<=18'h22834;
					11'h0365: dataout<=18'h0c6dc;
					11'h0366: dataout<=18'h06571;
					11'h0367: dataout<=18'h1f5d8;
					11'h0368: dataout<=18'h22a4d;
					11'h0369: dataout<=18'h0cbc5;
					11'h036a: dataout<=18'h0680e;
					11'h036b: dataout<=18'h1f54f;
					11'h036c: dataout<=18'h22c74;
					11'h036d: dataout<=18'h0d0a8;
					11'h036e: dataout<=18'h06aab;
					11'h036f: dataout<=18'h1f4c2;
					11'h0370: dataout<=18'h22ea7;
					11'h0371: dataout<=18'h0d585;
					11'h0372: dataout<=18'h06d47;
					11'h0373: dataout<=18'h1f432;
					11'h0374: dataout<=18'h230e8;
					11'h0375: dataout<=18'h0da5c;
					11'h0376: dataout<=18'h06fe2;
					11'h0377: dataout<=18'h1f39f;
					11'h0378: dataout<=18'h23335;
					11'h0379: dataout<=18'h0df2e;
					11'h037a: dataout<=18'h0727d;
					11'h037b: dataout<=18'h1f308;
					11'h037c: dataout<=18'h23590;
					11'h037d: dataout<=18'h0e3f9;
					11'h037e: dataout<=18'h07516;
					11'h037f: dataout<=18'h1f26d;
					11'h0380: dataout<=18'h237f7;
					11'h0381: dataout<=18'h0e8bd;
					11'h0382: dataout<=18'h077af;
					11'h0383: dataout<=18'h1f1cf;
					11'h0384: dataout<=18'h23a6a;
					11'h0385: dataout<=18'h0ed7b;
					11'h0386: dataout<=18'h07a47;
					11'h0387: dataout<=18'h1f12d;
					11'h0388: dataout<=18'h23cea;
					11'h0389: dataout<=18'h0f233;
					11'h038a: dataout<=18'h07cdf;
					11'h038b: dataout<=18'h1f088;
					11'h038c: dataout<=18'h23f77;
					11'h038d: dataout<=18'h0f6e4;
					11'h038e: dataout<=18'h07f75;
					11'h038f: dataout<=18'h1efe0;
					11'h0390: dataout<=18'h24211;
					11'h0391: dataout<=18'h0fb8e;
					11'h0392: dataout<=18'h0820a;
					11'h0393: dataout<=18'h1ef34;
					11'h0394: dataout<=18'h244b6;
					11'h0395: dataout<=18'h10031;
					11'h0396: dataout<=18'h0849f;
					11'h0397: dataout<=18'h1ee85;
					11'h0398: dataout<=18'h24769;
					11'h0399: dataout<=18'h104cd;
					11'h039a: dataout<=18'h08733;
					11'h039b: dataout<=18'h1edd2;
					11'h039c: dataout<=18'h24a27;
					11'h039d: dataout<=18'h10961;
					11'h039e: dataout<=18'h089c5;
					11'h039f: dataout<=18'h1ed1c;
					11'h03a0: dataout<=18'h24cf1;
					11'h03a1: dataout<=18'h10dee;
					11'h03a2: dataout<=18'h08c57;
					11'h03a3: dataout<=18'h1ec62;
					11'h03a4: dataout<=18'h24fc8;
					11'h03a5: dataout<=18'h11274;
					11'h03a6: dataout<=18'h08ee8;
					11'h03a7: dataout<=18'h1eba5;
					11'h03a8: dataout<=18'h252ab;
					11'h03a9: dataout<=18'h116f2;
					11'h03aa: dataout<=18'h09177;
					11'h03ab: dataout<=18'h1eae5;
					11'h03ac: dataout<=18'h25599;
					11'h03ad: dataout<=18'h11b68;
					11'h03ae: dataout<=18'h09406;
					11'h03af: dataout<=18'h1ea21;
					11'h03b0: dataout<=18'h25894;
					11'h03b1: dataout<=18'h11fd7;
					11'h03b2: dataout<=18'h09694;
					11'h03b3: dataout<=18'h1e95a;
					11'h03b4: dataout<=18'h25b9a;
					11'h03b5: dataout<=18'h1243d;
					11'h03b6: dataout<=18'h09921;
					11'h03b7: dataout<=18'h1e88f;
					11'h03b8: dataout<=18'h25eac;
					11'h03b9: dataout<=18'h1289b;
					11'h03ba: dataout<=18'h09bac;
					11'h03bb: dataout<=18'h1e7c1;
					11'h03bc: dataout<=18'h261ca;
					11'h03bd: dataout<=18'h12cf1;
					11'h03be: dataout<=18'h09e37;
					11'h03bf: dataout<=18'h1e6ef;
					11'h03c0: dataout<=18'h264f3;
					11'h03c1: dataout<=18'h1313f;
					11'h03c2: dataout<=18'h0a0c0;
					11'h03c3: dataout<=18'h1e61b;
					11'h03c4: dataout<=18'h26828;
					11'h03c5: dataout<=18'h13584;
					11'h03c6: dataout<=18'h0a348;
					11'h03c7: dataout<=18'h1e542;
					11'h03c8: dataout<=18'h26b68;
					11'h03c9: dataout<=18'h139c0;
					11'h03ca: dataout<=18'h0a5d0;
					11'h03cb: dataout<=18'h1e467;
					11'h03cc: dataout<=18'h26eb3;
					11'h03cd: dataout<=18'h13df4;
					11'h03ce: dataout<=18'h0a856;
					11'h03cf: dataout<=18'h1e388;
					11'h03d0: dataout<=18'h27209;
					11'h03d1: dataout<=18'h1421f;
					11'h03d2: dataout<=18'h0aada;
					11'h03d3: dataout<=18'h1e2a5;
					11'h03d4: dataout<=18'h2756b;
					11'h03d5: dataout<=18'h14641;
					11'h03d6: dataout<=18'h0ad5e;
					11'h03d7: dataout<=18'h1e1c0;
					11'h03d8: dataout<=18'h278d7;
					11'h03d9: dataout<=18'h14a5a;
					11'h03da: dataout<=18'h0afe0;
					11'h03db: dataout<=18'h1e0d6;
					11'h03dc: dataout<=18'h27c4e;
					11'h03dd: dataout<=18'h14e69;
					11'h03de: dataout<=18'h0b262;
					11'h03df: dataout<=18'h1dfea;
					11'h03e0: dataout<=18'h27fd1;
					11'h03e1: dataout<=18'h15270;
					11'h03e2: dataout<=18'h0b4e2;
					11'h03e3: dataout<=18'h1defa;
					11'h03e4: dataout<=18'h2835d;
					11'h03e5: dataout<=18'h1566c;
					11'h03e6: dataout<=18'h0b760;
					11'h03e7: dataout<=18'h1de07;
					11'h03e8: dataout<=18'h286f5;
					11'h03e9: dataout<=18'h15a60;
					11'h03ea: dataout<=18'h0b9de;
					11'h03eb: dataout<=18'h1dd11;
					11'h03ec: dataout<=18'h28a97;
					11'h03ed: dataout<=18'h15e4a;
					11'h03ee: dataout<=18'h0bc5a;
					11'h03ef: dataout<=18'h1dc17;
					11'h03f0: dataout<=18'h28e43;
					11'h03f1: dataout<=18'h16229;
					11'h03f2: dataout<=18'h0bed5;
					11'h03f3: dataout<=18'h1db1a;
					11'h03f4: dataout<=18'h291fa;
					11'h03f5: dataout<=18'h16600;
					11'h03f6: dataout<=18'h0c14e;
					11'h03f7: dataout<=18'h1da19;
					11'h03f8: dataout<=18'h295ba;
					11'h03f9: dataout<=18'h169cc;
					11'h03fa: dataout<=18'h0c3c6;
					11'h03fb: dataout<=18'h1d916;
					11'h03fc: dataout<=18'h29985;
					11'h03fd: dataout<=18'h16d8e;
					11'h03fe: dataout<=18'h0c63d;
					11'h03ff: dataout<=18'h1d80f;
					11'h0400: dataout<=18'h29d5a;
					11'h0401: dataout<=18'h17146;
					11'h0402: dataout<=18'h0c8b3;
					11'h0403: dataout<=18'h1d705;
					11'h0404: dataout<=18'h2a139;
					11'h0405: dataout<=18'h174f3;
					11'h0406: dataout<=18'h0cb27;
					11'h0407: dataout<=18'h1d5f7;
					11'h0408: dataout<=18'h2a521;
					11'h0409: dataout<=18'h17897;
					11'h040a: dataout<=18'h0cd99;
					11'h040b: dataout<=18'h1d4e6;
					11'h040c: dataout<=18'h2a914;
					11'h040d: dataout<=18'h17c2f;
					11'h040e: dataout<=18'h0d00a;
					11'h040f: dataout<=18'h1d3d2;
					11'h0410: dataout<=18'h2ad0f;
					11'h0411: dataout<=18'h17fbe;
					11'h0412: dataout<=18'h0d27a;
					11'h0413: dataout<=18'h1d2bb;
					11'h0414: dataout<=18'h2b114;
					11'h0415: dataout<=18'h18341;
					11'h0416: dataout<=18'h0d4e8;
					11'h0417: dataout<=18'h1d1a0;
					11'h0418: dataout<=18'h2b523;
					11'h0419: dataout<=18'h186ba;
					11'h041a: dataout<=18'h0d755;
					11'h041b: dataout<=18'h1d082;
					11'h041c: dataout<=18'h2b93b;
					11'h041d: dataout<=18'h18a28;
					11'h041e: dataout<=18'h0d9c0;
					11'h041f: dataout<=18'h1cf61;
					11'h0420: dataout<=18'h2bd5b;
					11'h0421: dataout<=18'h18d8a;
					11'h0422: dataout<=18'h0dc2a;
					11'h0423: dataout<=18'h1ce3d;
					11'h0424: dataout<=18'h2c185;
					11'h0425: dataout<=18'h190e2;
					11'h0426: dataout<=18'h0de92;
					11'h0427: dataout<=18'h1cd16;
					11'h0428: dataout<=18'h2c5b8;
					11'h0429: dataout<=18'h1942f;
					11'h042a: dataout<=18'h0e0f9;
					11'h042b: dataout<=18'h1cbeb;
					11'h042c: dataout<=18'h2c9f3;
					11'h042d: dataout<=18'h19770;
					11'h042e: dataout<=18'h0e35e;
					11'h042f: dataout<=18'h1cabd;
					11'h0430: dataout<=18'h2ce37;
					11'h0431: dataout<=18'h19aa6;
					11'h0432: dataout<=18'h0e5c2;
					11'h0433: dataout<=18'h1c98c;
					11'h0434: dataout<=18'h2d284;
					11'h0435: dataout<=18'h19dd1;
					11'h0436: dataout<=18'h0e824;
					11'h0437: dataout<=18'h1c858;
					11'h0438: dataout<=18'h2d6d8;
					11'h0439: dataout<=18'h1a0f0;
					11'h043a: dataout<=18'h0ea84;
					11'h043b: dataout<=18'h1c720;
					11'h043c: dataout<=18'h2db36;
					11'h043d: dataout<=18'h1a403;
					11'h043e: dataout<=18'h0ece3;
					11'h043f: dataout<=18'h1c5e6;
					11'h0440: dataout<=18'h2df9b;
					11'h0441: dataout<=18'h1a70b;
					11'h0442: dataout<=18'h0ef40;
					11'h0443: dataout<=18'h1c4a8;
					11'h0444: dataout<=18'h2e408;
					11'h0445: dataout<=18'h1aa07;
					11'h0446: dataout<=18'h0f19b;
					11'h0447: dataout<=18'h1c367;
					11'h0448: dataout<=18'h2e87e;
					11'h0449: dataout<=18'h1acf7;
					11'h044a: dataout<=18'h0f3f5;
					11'h044b: dataout<=18'h1c223;
					11'h044c: dataout<=18'h2ecfb;
					11'h044d: dataout<=18'h1afdb;
					11'h044e: dataout<=18'h0f64d;
					11'h044f: dataout<=18'h1c0dc;
					11'h0450: dataout<=18'h2f17f;
					11'h0451: dataout<=18'h1b2b4;
					11'h0452: dataout<=18'h0f8a3;
					11'h0453: dataout<=18'h1bf91;
					11'h0454: dataout<=18'h2f60c;
					11'h0455: dataout<=18'h1b580;
					11'h0456: dataout<=18'h0faf8;
					11'h0457: dataout<=18'h1be44;
					11'h0458: dataout<=18'h2fa9f;
					11'h0459: dataout<=18'h1b840;
					11'h045a: dataout<=18'h0fd4a;
					11'h045b: dataout<=18'h1bcf3;
					11'h045c: dataout<=18'h2ff3a;
					11'h045d: dataout<=18'h1baf3;
					11'h045e: dataout<=18'h0ff9c;
					11'h045f: dataout<=18'h1bba0;
					11'h0460: dataout<=18'h303dc;
					11'h0461: dataout<=18'h1bd9b;
					11'h0462: dataout<=18'h101eb;
					11'h0463: dataout<=18'h1ba49;
					11'h0464: dataout<=18'h30885;
					11'h0465: dataout<=18'h1c035;
					11'h0466: dataout<=18'h10438;
					11'h0467: dataout<=18'h1b8ef;
					11'h0468: dataout<=18'h30d35;
					11'h0469: dataout<=18'h1c2c4;
					11'h046a: dataout<=18'h10684;
					11'h046b: dataout<=18'h1b792;
					11'h046c: dataout<=18'h311ec;
					11'h046d: dataout<=18'h1c546;
					11'h046e: dataout<=18'h108ce;
					11'h046f: dataout<=18'h1b632;
					11'h0470: dataout<=18'h316a9;
					11'h0471: dataout<=18'h1c7bb;
					11'h0472: dataout<=18'h10b16;
					11'h0473: dataout<=18'h1b4cf;
					11'h0474: dataout<=18'h31b6d;
					11'h0475: dataout<=18'h1ca24;
					11'h0476: dataout<=18'h10d5c;
					11'h0477: dataout<=18'h1b369;
					11'h0478: dataout<=18'h32037;
					11'h0479: dataout<=18'h1cc7f;
					11'h047a: dataout<=18'h10fa0;
					11'h047b: dataout<=18'h1b200;
					11'h047c: dataout<=18'h32508;
					11'h047d: dataout<=18'h1cece;
					11'h047e: dataout<=18'h111e2;
					11'h047f: dataout<=18'h1b094;
					11'h0480: dataout<=18'h329de;
					11'h0481: dataout<=18'h1d111;
					11'h0482: dataout<=18'h11423;
					11'h0483: dataout<=18'h1af25;
					11'h0484: dataout<=18'h32ebb;
					11'h0485: dataout<=18'h1d346;
					11'h0486: dataout<=18'h11661;
					11'h0487: dataout<=18'h1adb3;
					11'h0488: dataout<=18'h3339d;
					11'h0489: dataout<=18'h1d56e;
					11'h048a: dataout<=18'h1189e;
					11'h048b: dataout<=18'h1ac3e;
					11'h048c: dataout<=18'h33885;
					11'h048d: dataout<=18'h1d789;
					11'h048e: dataout<=18'h11ad9;
					11'h048f: dataout<=18'h1aac6;
					11'h0490: dataout<=18'h33d73;
					11'h0491: dataout<=18'h1d997;
					11'h0492: dataout<=18'h11d11;
					11'h0493: dataout<=18'h1a94b;
					11'h0494: dataout<=18'h34266;
					11'h0495: dataout<=18'h1db98;
					11'h0496: dataout<=18'h11f48;
					11'h0497: dataout<=18'h1a7cd;
					11'h0498: dataout<=18'h3475e;
					11'h0499: dataout<=18'h1dd8b;
					11'h049a: dataout<=18'h1217d;
					11'h049b: dataout<=18'h1a64c;
					11'h049c: dataout<=18'h34c5c;
					11'h049d: dataout<=18'h1df72;
					11'h049e: dataout<=18'h123af;
					11'h049f: dataout<=18'h1a4c8;
					11'h04a0: dataout<=18'h3515e;
					11'h04a1: dataout<=18'h1e14a;
					11'h04a2: dataout<=18'h125e0;
					11'h04a3: dataout<=18'h1a341;
					11'h04a4: dataout<=18'h35665;
					11'h04a5: dataout<=18'h1e316;
					11'h04a6: dataout<=18'h1280f;
					11'h04a7: dataout<=18'h1a1b8;
					11'h04a8: dataout<=18'h35b71;
					11'h04a9: dataout<=18'h1e4d4;
					11'h04aa: dataout<=18'h12a3b;
					11'h04ab: dataout<=18'h1a02b;
					11'h04ac: dataout<=18'h36082;
					11'h04ad: dataout<=18'h1e685;
					11'h04ae: dataout<=18'h12c66;
					11'h04af: dataout<=18'h19e9b;
					11'h04b0: dataout<=18'h36597;
					11'h04b1: dataout<=18'h1e828;
					11'h04b2: dataout<=18'h12e8e;
					11'h04b3: dataout<=18'h19d09;
					11'h04b4: dataout<=18'h36ab0;
					11'h04b5: dataout<=18'h1e9bd;
					11'h04b6: dataout<=18'h130b4;
					11'h04b7: dataout<=18'h19b74;
					11'h04b8: dataout<=18'h36fce;
					11'h04b9: dataout<=18'h1eb45;
					11'h04ba: dataout<=18'h132d8;
					11'h04bb: dataout<=18'h199db;
					11'h04bc: dataout<=18'h374ef;
					11'h04bd: dataout<=18'h1ecbf;
					11'h04be: dataout<=18'h134fa;
					11'h04bf: dataout<=18'h19840;
					11'h04c0: dataout<=18'h37a14;
					11'h04c1: dataout<=18'h1ee2b;
					11'h04c2: dataout<=18'h1371a;
					11'h04c3: dataout<=18'h196a3;
					11'h04c4: dataout<=18'h37f3d;
					11'h04c5: dataout<=18'h1ef8a;
					11'h04c6: dataout<=18'h13938;
					11'h04c7: dataout<=18'h19502;
					11'h04c8: dataout<=18'h3846a;
					11'h04c9: dataout<=18'h1f0db;
					11'h04ca: dataout<=18'h13b54;
					11'h04cb: dataout<=18'h1935e;
					11'h04cc: dataout<=18'h3899a;
					11'h04cd: dataout<=18'h1f21e;
					11'h04ce: dataout<=18'h13d6d;
					11'h04cf: dataout<=18'h191b8;
					11'h04d0: dataout<=18'h38ece;
					11'h04d1: dataout<=18'h1f353;
					11'h04d2: dataout<=18'h13f84;
					11'h04d3: dataout<=18'h1900f;
					11'h04d4: dataout<=18'h39404;
					11'h04d5: dataout<=18'h1f47a;
					11'h04d6: dataout<=18'h14199;
					11'h04d7: dataout<=18'h18e63;
					11'h04d8: dataout<=18'h3993e;
					11'h04d9: dataout<=18'h1f593;
					11'h04da: dataout<=18'h143ab;
					11'h04db: dataout<=18'h18cb5;
					11'h04dc: dataout<=18'h39e7a;
					11'h04dd: dataout<=18'h1f69f;
					11'h04de: dataout<=18'h145bc;
					11'h04df: dataout<=18'h18b03;
					11'h04e0: dataout<=18'h3a3b9;
					11'h04e1: dataout<=18'h1f79c;
					11'h04e2: dataout<=18'h147ca;
					11'h04e3: dataout<=18'h1894f;
					11'h04e4: dataout<=18'h3a8fb;
					11'h04e5: dataout<=18'h1f88b;
					11'h04e6: dataout<=18'h149d6;
					11'h04e7: dataout<=18'h18798;
					11'h04e8: dataout<=18'h3ae3f;
					11'h04e9: dataout<=18'h1f96d;
					11'h04ea: dataout<=18'h14bdf;
					11'h04eb: dataout<=18'h185de;
					11'h04ec: dataout<=18'h3b386;
					11'h04ed: dataout<=18'h1fa40;
					11'h04ee: dataout<=18'h14de7;
					11'h04ef: dataout<=18'h18422;
					11'h04f0: dataout<=18'h3b8ce;
					11'h04f1: dataout<=18'h1fb05;
					11'h04f2: dataout<=18'h14fec;
					11'h04f3: dataout<=18'h18263;
					11'h04f4: dataout<=18'h3be19;
					11'h04f5: dataout<=18'h1fbbc;
					11'h04f6: dataout<=18'h151ee;
					11'h04f7: dataout<=18'h180a1;
					11'h04f8: dataout<=18'h3c365;
					11'h04f9: dataout<=18'h1fc65;
					11'h04fa: dataout<=18'h153ee;
					11'h04fb: dataout<=18'h17edd;
					11'h04fc: dataout<=18'h3c8b3;
					11'h04fd: dataout<=18'h1fd00;
					11'h04fe: dataout<=18'h155ec;
					11'h04ff: dataout<=18'h17d16;
					11'h0500: dataout<=18'h3ce03;
					11'h0501: dataout<=18'h1fd8c;
					11'h0502: dataout<=18'h157e8;
					11'h0503: dataout<=18'h17b4c;
					11'h0504: dataout<=18'h3d354;
					11'h0505: dataout<=18'h1fe0b;
					11'h0506: dataout<=18'h159e1;
					11'h0507: dataout<=18'h17980;
					11'h0508: dataout<=18'h3d8a6;
					11'h0509: dataout<=18'h1fe7b;
					11'h050a: dataout<=18'h15bd8;
					11'h050b: dataout<=18'h177b1;
					11'h050c: dataout<=18'h3ddf9;
					11'h050d: dataout<=18'h1fedd;
					11'h050e: dataout<=18'h15dcc;
					11'h050f: dataout<=18'h175df;
					11'h0510: dataout<=18'h3e34d;
					11'h0511: dataout<=18'h1ff30;
					11'h0512: dataout<=18'h15fbe;
					11'h0513: dataout<=18'h1740b;
					11'h0514: dataout<=18'h3e8a2;
					11'h0515: dataout<=18'h1ff76;
					11'h0516: dataout<=18'h161ad;
					11'h0517: dataout<=18'h17234;
					11'h0518: dataout<=18'h3edf8;
					11'h0519: dataout<=18'h1ffad;
					11'h051a: dataout<=18'h1639a;
					11'h051b: dataout<=18'h1705b;
					11'h051c: dataout<=18'h3f34e;
					11'h051d: dataout<=18'h1ffd6;
					11'h051e: dataout<=18'h16584;
					11'h051f: dataout<=18'h16e7f;
					11'h0520: dataout<=18'h3f8a5;
					11'h0521: dataout<=18'h1fff1;
					11'h0522: dataout<=18'h1676c;
					11'h0523: dataout<=18'h16ca0;
					11'h0524: dataout<=18'h3fdfc;
					11'h0525: dataout<=18'h1fffd;
					11'h0526: dataout<=18'h16952;
					11'h0527: dataout<=18'h16abf;
					11'h0528: dataout<=18'h00351;
					11'h0529: dataout<=18'h1fffc;
					11'h052a: dataout<=18'h16b35;
					11'h052b: dataout<=18'h168dc;
					11'h052c: dataout<=18'h008a8;
					11'h052d: dataout<=18'h1ffec;
					11'h052e: dataout<=18'h16d15;
					11'h052f: dataout<=18'h166f6;
					11'h0530: dataout<=18'h00dff;
					11'h0531: dataout<=18'h1ffce;
					11'h0532: dataout<=18'h16ef3;
					11'h0533: dataout<=18'h1650d;
					11'h0534: dataout<=18'h01355;
					11'h0535: dataout<=18'h1ffa1;
					11'h0536: dataout<=18'h170ce;
					11'h0537: dataout<=18'h16322;
					11'h0538: dataout<=18'h018aa;
					11'h0539: dataout<=18'h1ff66;
					11'h053a: dataout<=18'h172a7;
					11'h053b: dataout<=18'h16135;
					11'h053c: dataout<=18'h01dff;
					11'h053d: dataout<=18'h1ff1d;
					11'h053e: dataout<=18'h1747d;
					11'h053f: dataout<=18'h15f45;
					11'h0540: dataout<=18'h02353;
					11'h0541: dataout<=18'h1fec6;
					11'h0542: dataout<=18'h17651;
					11'h0543: dataout<=18'h15d52;
					11'h0544: dataout<=18'h028a6;
					11'h0545: dataout<=18'h1fe61;
					11'h0546: dataout<=18'h17822;
					11'h0547: dataout<=18'h15b5d;
					11'h0548: dataout<=18'h02df8;
					11'h0549: dataout<=18'h1fded;
					11'h054a: dataout<=18'h179f0;
					11'h054b: dataout<=18'h15966;
					11'h054c: dataout<=18'h03349;
					11'h054d: dataout<=18'h1fd6b;
					11'h054e: dataout<=18'h17bbc;
					11'h054f: dataout<=18'h1576c;
					11'h0550: dataout<=18'h03898;
					11'h0551: dataout<=18'h1fcdb;
					11'h0552: dataout<=18'h17d85;
					11'h0553: dataout<=18'h15570;
					11'h0554: dataout<=18'h03de6;
					11'h0555: dataout<=18'h1fc3d;
					11'h0556: dataout<=18'h17f4b;
					11'h0557: dataout<=18'h15372;
					11'h0558: dataout<=18'h04332;
					11'h0559: dataout<=18'h1fb91;
					11'h055a: dataout<=18'h1810f;
					11'h055b: dataout<=18'h15171;
					11'h055c: dataout<=18'h0487c;
					11'h055d: dataout<=18'h1fad6;
					11'h055e: dataout<=18'h182d0;
					11'h055f: dataout<=18'h14f6e;
					11'h0560: dataout<=18'h04dc4;
					11'h0561: dataout<=18'h1fa0e;
					11'h0562: dataout<=18'h1848f;
					11'h0563: dataout<=18'h14d68;
					11'h0564: dataout<=18'h0530a;
					11'h0565: dataout<=18'h1f937;
					11'h0566: dataout<=18'h1864a;
					11'h0567: dataout<=18'h14b61;
					11'h0568: dataout<=18'h0584d;
					11'h0569: dataout<=18'h1f852;
					11'h056a: dataout<=18'h18803;
					11'h056b: dataout<=18'h14956;
					11'h056c: dataout<=18'h05d8e;
					11'h056d: dataout<=18'h1f760;
					11'h056e: dataout<=18'h189b9;
					11'h056f: dataout<=18'h1474a;
					11'h0570: dataout<=18'h062cd;
					11'h0571: dataout<=18'h1f65f;
					11'h0572: dataout<=18'h18b6d;
					11'h0573: dataout<=18'h1453b;
					11'h0574: dataout<=18'h06808;
					11'h0575: dataout<=18'h1f550;
					11'h0576: dataout<=18'h18d1e;
					11'h0577: dataout<=18'h1432a;
					11'h0578: dataout<=18'h06d41;
					11'h0579: dataout<=18'h1f433;
					11'h057a: dataout<=18'h18ecc;
					11'h057b: dataout<=18'h14117;
					11'h057c: dataout<=18'h07277;
					11'h057d: dataout<=18'h1f309;
					11'h057e: dataout<=18'h19077;
					11'h057f: dataout<=18'h13f02;
					11'h0580: dataout<=18'h077aa;
					11'h0581: dataout<=18'h1f1d0;
					11'h0582: dataout<=18'h1921f;
					11'h0583: dataout<=18'h13cea;
					11'h0584: dataout<=18'h07cd9;
					11'h0585: dataout<=18'h1f08a;
					11'h0586: dataout<=18'h193c5;
					11'h0587: dataout<=18'h13ad0;
					11'h0588: dataout<=18'h08205;
					11'h0589: dataout<=18'h1ef36;
					11'h058a: dataout<=18'h19568;
					11'h058b: dataout<=18'h138b4;
					11'h058c: dataout<=18'h0872d;
					11'h058d: dataout<=18'h1edd4;
					11'h058e: dataout<=18'h19708;
					11'h058f: dataout<=18'h13696;
					11'h0590: dataout<=18'h08c51;
					11'h0591: dataout<=18'h1ec64;
					11'h0592: dataout<=18'h198a5;
					11'h0593: dataout<=18'h13476;
					11'h0594: dataout<=18'h09172;
					11'h0595: dataout<=18'h1eae7;
					11'h0596: dataout<=18'h19a3f;
					11'h0597: dataout<=18'h13253;
					11'h0598: dataout<=18'h0968e;
					11'h0599: dataout<=18'h1e95b;
					11'h059a: dataout<=18'h19bd7;
					11'h059b: dataout<=18'h1302e;
					11'h059c: dataout<=18'h09ba7;
					11'h059d: dataout<=18'h1e7c3;
					11'h059e: dataout<=18'h19d6b;
					11'h059f: dataout<=18'h12e08;
					11'h05a0: dataout<=18'h0a0bb;
					11'h05a1: dataout<=18'h1e61c;
					11'h05a2: dataout<=18'h19efd;
					11'h05a3: dataout<=18'h12bdf;
					11'h05a4: dataout<=18'h0a5ca;
					11'h05a5: dataout<=18'h1e469;
					11'h05a6: dataout<=18'h1a08c;
					11'h05a7: dataout<=18'h129b4;
					11'h05a8: dataout<=18'h0aad5;
					11'h05a9: dataout<=18'h1e2a7;
					11'h05aa: dataout<=18'h1a218;
					11'h05ab: dataout<=18'h12787;
					11'h05ac: dataout<=18'h0afdb;
					11'h05ad: dataout<=18'h1e0d8;
					11'h05ae: dataout<=18'h1a3a1;
					11'h05af: dataout<=18'h12558;
					11'h05b0: dataout<=18'h0b4dc;
					11'h05b1: dataout<=18'h1defc;
					11'h05b2: dataout<=18'h1a527;
					11'h05b3: dataout<=18'h12326;
					11'h05b4: dataout<=18'h0b9d8;
					11'h05b5: dataout<=18'h1dd13;
					11'h05b6: dataout<=18'h1a6aa;
					11'h05b7: dataout<=18'h120f3;
					11'h05b8: dataout<=18'h0becf;
					11'h05b9: dataout<=18'h1db1c;
					11'h05ba: dataout<=18'h1a82a;
					11'h05bb: dataout<=18'h11ebe;
					11'h05bc: dataout<=18'h0c3c1;
					11'h05bd: dataout<=18'h1d918;
					11'h05be: dataout<=18'h1a9a7;
					11'h05bf: dataout<=18'h11c87;
					11'h05c0: dataout<=18'h0c8ad;
					11'h05c1: dataout<=18'h1d707;
					11'h05c2: dataout<=18'h1ab22;
					11'h05c3: dataout<=18'h11a4e;
					11'h05c4: dataout<=18'h0cd94;
					11'h05c5: dataout<=18'h1d4e9;
					11'h05c6: dataout<=18'h1ac99;
					11'h05c7: dataout<=18'h11813;
					11'h05c8: dataout<=18'h0d275;
					11'h05c9: dataout<=18'h1d2bd;
					11'h05ca: dataout<=18'h1ae0d;
					11'h05cb: dataout<=18'h115d6;
					11'h05cc: dataout<=18'h0d750;
					11'h05cd: dataout<=18'h1d085;
					11'h05ce: dataout<=18'h1af7f;
					11'h05cf: dataout<=18'h11397;
					11'h05d0: dataout<=18'h0dc25;
					11'h05d1: dataout<=18'h1ce40;
					11'h05d2: dataout<=18'h1b0ed;
					11'h05d3: dataout<=18'h11156;
					11'h05d4: dataout<=18'h0e0f4;
					11'h05d5: dataout<=18'h1cbed;
					11'h05d6: dataout<=18'h1b259;
					11'h05d7: dataout<=18'h10f13;
					11'h05d8: dataout<=18'h0e5bd;
					11'h05d9: dataout<=18'h1c98f;
					11'h05da: dataout<=18'h1b3c1;
					11'h05db: dataout<=18'h10cce;
					11'h05dc: dataout<=18'h0ea7f;
					11'h05dd: dataout<=18'h1c723;
					11'h05de: dataout<=18'h1b526;
					11'h05df: dataout<=18'h10a88;
					11'h05e0: dataout<=18'h0ef3b;
					11'h05e1: dataout<=18'h1c4ab;
					11'h05e2: dataout<=18'h1b688;
					11'h05e3: dataout<=18'h1083f;
					11'h05e4: dataout<=18'h0f3f0;
					11'h05e5: dataout<=18'h1c226;
					11'h05e6: dataout<=18'h1b7e8;
					11'h05e7: dataout<=18'h105f5;
					11'h05e8: dataout<=18'h0f89e;
					11'h05e9: dataout<=18'h1bf94;
					11'h05ea: dataout<=18'h1b944;
					11'h05eb: dataout<=18'h103a9;
					11'h05ec: dataout<=18'h0fd45;
					11'h05ed: dataout<=18'h1bcf6;
					11'h05ee: dataout<=18'h1ba9d;
					11'h05ef: dataout<=18'h1015b;
					11'h05f0: dataout<=18'h101e6;
					11'h05f1: dataout<=18'h1ba4c;
					11'h05f2: dataout<=18'h1bbf3;
					11'h05f3: dataout<=18'h0ff0b;
					11'h05f4: dataout<=18'h1067f;
					11'h05f5: dataout<=18'h1b795;
					11'h05f6: dataout<=18'h1bd46;
					11'h05f7: dataout<=18'h0fcba;
					11'h05f8: dataout<=18'h10b11;
					11'h05f9: dataout<=18'h1b4d2;
					11'h05fa: dataout<=18'h1be95;
					11'h05fb: dataout<=18'h0fa66;
					11'h05fc: dataout<=18'h10f9b;
					11'h05fd: dataout<=18'h1b203;
					11'h05fe: dataout<=18'h1bfe2;
					11'h05ff: dataout<=18'h0f811;
					11'h0600: dataout<=18'h1141e;
					11'h0601: dataout<=18'h1af28;
					11'h0602: dataout<=18'h1c12c;
					11'h0603: dataout<=18'h0f5bb;
					11'h0604: dataout<=18'h11899;
					11'h0605: dataout<=18'h1ac41;
					11'h0606: dataout<=18'h1c272;
					11'h0607: dataout<=18'h0f362;
					11'h0608: dataout<=18'h11d0d;
					11'h0609: dataout<=18'h1a94e;
					11'h060a: dataout<=18'h1c3b5;
					11'h060b: dataout<=18'h0f108;
					11'h060c: dataout<=18'h12178;
					11'h060d: dataout<=18'h1a64f;
					11'h060e: dataout<=18'h1c4f6;
					11'h060f: dataout<=18'h0eeac;
					11'h0610: dataout<=18'h125db;
					11'h0611: dataout<=18'h1a345;
					11'h0612: dataout<=18'h1c633;
					11'h0613: dataout<=18'h0ec4f;
					11'h0614: dataout<=18'h12a37;
					11'h0615: dataout<=18'h1a02e;
					11'h0616: dataout<=18'h1c76c;
					11'h0617: dataout<=18'h0e9f0;
					11'h0618: dataout<=18'h12e89;
					11'h0619: dataout<=18'h19d0c;
					11'h061a: dataout<=18'h1c8a3;
					11'h061b: dataout<=18'h0e78f;
					11'h061c: dataout<=18'h132d4;
					11'h061d: dataout<=18'h199df;
					11'h061e: dataout<=18'h1c9d7;
					11'h061f: dataout<=18'h0e52d;
					11'h0620: dataout<=18'h13716;
					11'h0621: dataout<=18'h196a6;
					11'h0622: dataout<=18'h1cb07;
					11'h0623: dataout<=18'h0e2c9;
					11'h0624: dataout<=18'h13b4f;
					11'h0625: dataout<=18'h19362;
					11'h0626: dataout<=18'h1cc34;
					11'h0627: dataout<=18'h0e063;
					11'h0628: dataout<=18'h13f7f;
					11'h0629: dataout<=18'h19013;
					11'h062a: dataout<=18'h1cd5e;
					11'h062b: dataout<=18'h0ddfc;
					11'h062c: dataout<=18'h143a7;
					11'h062d: dataout<=18'h18cb8;
					11'h062e: dataout<=18'h1ce85;
					11'h062f: dataout<=18'h0db94;
					11'h0630: dataout<=18'h147c6;
					11'h0631: dataout<=18'h18953;
					11'h0632: dataout<=18'h1cfa8;
					11'h0633: dataout<=18'h0d92a;
					11'h0634: dataout<=18'h14bdb;
					11'h0635: dataout<=18'h185e2;
					11'h0636: dataout<=18'h1d0c8;
					11'h0637: dataout<=18'h0d6be;
					11'h0638: dataout<=18'h14fe7;
					11'h0639: dataout<=18'h18267;
					11'h063a: dataout<=18'h1d1e5;
					11'h063b: dataout<=18'h0d451;
					11'h063c: dataout<=18'h153ea;
					11'h063d: dataout<=18'h17ee1;
					11'h063e: dataout<=18'h1d2ff;
					11'h063f: dataout<=18'h0d1e2;
					11'h0640: dataout<=18'h157e3;
					11'h0641: dataout<=18'h17b50;
					11'h0642: dataout<=18'h1d416;
					11'h0643: dataout<=18'h0cf72;
					11'h0644: dataout<=18'h15bd3;
					11'h0645: dataout<=18'h177b5;
					11'h0646: dataout<=18'h1d529;
					11'h0647: dataout<=18'h0cd01;
					11'h0648: dataout<=18'h15fb9;
					11'h0649: dataout<=18'h1740f;
					11'h064a: dataout<=18'h1d639;
					11'h064b: dataout<=18'h0ca8e;
					11'h064c: dataout<=18'h16396;
					11'h064d: dataout<=18'h1705f;
					11'h064e: dataout<=18'h1d746;
					11'h064f: dataout<=18'h0c819;
					11'h0650: dataout<=18'h16768;
					11'h0651: dataout<=18'h16ca4;
					11'h0652: dataout<=18'h1d84f;
					11'h0653: dataout<=18'h0c5a4;
					11'h0654: dataout<=18'h16b31;
					11'h0655: dataout<=18'h168e0;
					11'h0656: dataout<=18'h1d955;
					11'h0657: dataout<=18'h0c32c;
					11'h0658: dataout<=18'h16eef;
					11'h0659: dataout<=18'h16511;
					11'h065a: dataout<=18'h1da58;
					11'h065b: dataout<=18'h0c0b4;
					11'h065c: dataout<=18'h172a3;
					11'h065d: dataout<=18'h16139;
					11'h065e: dataout<=18'h1db58;
					11'h065f: dataout<=18'h0be3a;
					11'h0660: dataout<=18'h1764d;
					11'h0661: dataout<=18'h15d56;
					11'h0662: dataout<=18'h1dc54;
					11'h0663: dataout<=18'h0bbbf;
					11'h0664: dataout<=18'h179ec;
					11'h0665: dataout<=18'h1596a;
					11'h0666: dataout<=18'h1dd4d;
					11'h0667: dataout<=18'h0b943;
					11'h0668: dataout<=18'h17d81;
					11'h0669: dataout<=18'h15575;
					11'h066a: dataout<=18'h1de43;
					11'h066b: dataout<=18'h0b6c5;
					11'h066c: dataout<=18'h1810b;
					11'h066d: dataout<=18'h15175;
					11'h066e: dataout<=18'h1df35;
					11'h066f: dataout<=18'h0b446;
					11'h0670: dataout<=18'h1848b;
					11'h0671: dataout<=18'h14d6d;
					11'h0672: dataout<=18'h1e024;
					11'h0673: dataout<=18'h0b1c6;
					11'h0674: dataout<=18'h18800;
					11'h0675: dataout<=18'h1495b;
					11'h0676: dataout<=18'h1e110;
					11'h0677: dataout<=18'h0af44;
					11'h0678: dataout<=18'h18b69;
					11'h0679: dataout<=18'h14540;
					11'h067a: dataout<=18'h1e1f8;
					11'h067b: dataout<=18'h0acc1;
					11'h067c: dataout<=18'h18ec8;
					11'h067d: dataout<=18'h1411c;
					11'h067e: dataout<=18'h1e2dd;
					11'h067f: dataout<=18'h0aa3d;
					11'h0680: dataout<=18'h1921c;
					11'h0681: dataout<=18'h13cef;
					11'h0682: dataout<=18'h1e3be;
					11'h0683: dataout<=18'h0a7b8;
					11'h0684: dataout<=18'h19564;
					11'h0685: dataout<=18'h138b9;
					11'h0686: dataout<=18'h1e49c;
					11'h0687: dataout<=18'h0a532;
					11'h0688: dataout<=18'h198a1;
					11'h0689: dataout<=18'h1347a;
					11'h068a: dataout<=18'h1e577;
					11'h068b: dataout<=18'h0a2aa;
					11'h068c: dataout<=18'h19bd3;
					11'h068d: dataout<=18'h13033;
					11'h068e: dataout<=18'h1e64f;
					11'h068f: dataout<=18'h0a022;
					11'h0690: dataout<=18'h19efa;
					11'h0691: dataout<=18'h12be3;
					11'h0692: dataout<=18'h1e723;
					11'h0693: dataout<=18'h09d98;
					11'h0694: dataout<=18'h1a214;
					11'h0695: dataout<=18'h1278b;
					11'h0696: dataout<=18'h1e7f3;
					11'h0697: dataout<=18'h09b0d;
					11'h0698: dataout<=18'h1a524;
					11'h0699: dataout<=18'h1232b;
					11'h069a: dataout<=18'h1e8c1;
					11'h069b: dataout<=18'h09882;
					11'h069c: dataout<=18'h1a827;
					11'h069d: dataout<=18'h11ec3;
					11'h069e: dataout<=18'h1e98b;
					11'h069f: dataout<=18'h095f5;
					11'h06a0: dataout<=18'h1ab1f;
					11'h06a1: dataout<=18'h11a53;
					11'h06a2: dataout<=18'h1ea51;
					11'h06a3: dataout<=18'h09367;
					11'h06a4: dataout<=18'h1ae0a;
					11'h06a5: dataout<=18'h115da;
					11'h06a6: dataout<=18'h1eb14;
					11'h06a7: dataout<=18'h090d8;
					11'h06a8: dataout<=18'h1b0ea;
					11'h06a9: dataout<=18'h1115b;
					11'h06aa: dataout<=18'h1ebd4;
					11'h06ab: dataout<=18'h08e48;
					11'h06ac: dataout<=18'h1b3be;
					11'h06ad: dataout<=18'h10cd3;
					11'h06ae: dataout<=18'h1ec90;
					11'h06af: dataout<=18'h08bb7;
					11'h06b0: dataout<=18'h1b685;
					11'h06b1: dataout<=18'h10844;
					11'h06b2: dataout<=18'h1ed49;
					11'h06b3: dataout<=18'h08925;
					11'h06b4: dataout<=18'h1b941;
					11'h06b5: dataout<=18'h103ae;
					11'h06b6: dataout<=18'h1edfe;
					11'h06b7: dataout<=18'h08692;
					11'h06b8: dataout<=18'h1bbf0;
					11'h06b9: dataout<=18'h0ff10;
					11'h06ba: dataout<=18'h1eeb0;
					11'h06bb: dataout<=18'h083fe;
					11'h06bc: dataout<=18'h1be93;
					11'h06bd: dataout<=18'h0fa6b;
					11'h06be: dataout<=18'h1ef5e;
					11'h06bf: dataout<=18'h08169;
					11'h06c0: dataout<=18'h1c129;
					11'h06c1: dataout<=18'h0f5c0;
					11'h06c2: dataout<=18'h1f009;
					11'h06c3: dataout<=18'h07ed4;
					11'h06c4: dataout<=18'h1c3b3;
					11'h06c5: dataout<=18'h0f10d;
					11'h06c6: dataout<=18'h1f0b1;
					11'h06c7: dataout<=18'h07c3d;
					11'h06c8: dataout<=18'h1c630;
					11'h06c9: dataout<=18'h0ec54;
					11'h06ca: dataout<=18'h1f155;
					11'h06cb: dataout<=18'h079a6;
					11'h06cc: dataout<=18'h1c8a1;
					11'h06cd: dataout<=18'h0e794;
					11'h06ce: dataout<=18'h1f1f6;
					11'h06cf: dataout<=18'h0770d;
					11'h06d0: dataout<=18'h1cb04;
					11'h06d1: dataout<=18'h0e2ce;
					11'h06d2: dataout<=18'h1f293;
					11'h06d3: dataout<=18'h07474;
					11'h06d4: dataout<=18'h1cd5b;
					11'h06d5: dataout<=18'h0de02;
					11'h06d6: dataout<=18'h1f32d;
					11'h06d7: dataout<=18'h071da;
					11'h06d8: dataout<=18'h1cfa6;
					11'h06d9: dataout<=18'h0d92f;
					11'h06da: dataout<=18'h1f3c3;
					11'h06db: dataout<=18'h06f40;
					11'h06dc: dataout<=18'h1d1e3;
					11'h06dd: dataout<=18'h0d456;
					11'h06de: dataout<=18'h1f456;
					11'h06df: dataout<=18'h06ca4;
					11'h06e0: dataout<=18'h1d413;
					11'h06e1: dataout<=18'h0cf77;
					11'h06e2: dataout<=18'h1f4e5;
					11'h06e3: dataout<=18'h06a08;
					11'h06e4: dataout<=18'h1d637;
					11'h06e5: dataout<=18'h0ca93;
					11'h06e6: dataout<=18'h1f571;
					11'h06e7: dataout<=18'h0676b;
					11'h06e8: dataout<=18'h1d84d;
					11'h06e9: dataout<=18'h0c5a9;
					11'h06ea: dataout<=18'h1f5f9;
					11'h06eb: dataout<=18'h064cd;
					11'h06ec: dataout<=18'h1da56;
					11'h06ed: dataout<=18'h0c0b9;
					11'h06ee: dataout<=18'h1f67e;
					11'h06ef: dataout<=18'h0622f;
					11'h06f0: dataout<=18'h1dc52;
					11'h06f1: dataout<=18'h0bbc4;
					11'h06f2: dataout<=18'h1f6ff;
					11'h06f3: dataout<=18'h05f90;
					11'h06f4: dataout<=18'h1de41;
					11'h06f5: dataout<=18'h0b6ca;
					11'h06f6: dataout<=18'h1f77d;
					11'h06f7: dataout<=18'h05cf0;
					11'h06f8: dataout<=18'h1e022;
					11'h06f9: dataout<=18'h0b1cb;
					11'h06fa: dataout<=18'h1f7f7;
					11'h06fb: dataout<=18'h05a50;
					11'h06fc: dataout<=18'h1e1f6;
					11'h06fd: dataout<=18'h0acc7;
					11'h06fe: dataout<=18'h1f86e;
					11'h06ff: dataout<=18'h057af;
					11'h0700: dataout<=18'h1e3bc;
					11'h0701: dataout<=18'h0a7be;
					11'h0702: dataout<=18'h1f8e1;
					11'h0703: dataout<=18'h0550d;
					11'h0704: dataout<=18'h1e575;
					11'h0705: dataout<=18'h0a2b0;
					11'h0706: dataout<=18'h1f951;
					11'h0707: dataout<=18'h0526b;
					11'h0708: dataout<=18'h1e721;
					11'h0709: dataout<=18'h09d9e;
					11'h070a: dataout<=18'h1f9bd;
					11'h070b: dataout<=18'h04fc8;
					11'h070c: dataout<=18'h1e8bf;
					11'h070d: dataout<=18'h09887;
					11'h070e: dataout<=18'h1fa26;
					11'h070f: dataout<=18'h04d25;
					11'h0710: dataout<=18'h1ea4f;
					11'h0711: dataout<=18'h0936c;
					11'h0712: dataout<=18'h1fa8b;
					11'h0713: dataout<=18'h04a81;
					11'h0714: dataout<=18'h1ebd2;
					11'h0715: dataout<=18'h08e4d;
					11'h0716: dataout<=18'h1faed;
					11'h0717: dataout<=18'h047dc;
					11'h0718: dataout<=18'h1ed47;
					11'h0719: dataout<=18'h0892a;
					11'h071a: dataout<=18'h1fb4b;
					11'h071b: dataout<=18'h04538;
					11'h071c: dataout<=18'h1eeae;
					11'h071d: dataout<=18'h08404;
					11'h071e: dataout<=18'h1fba6;
					11'h071f: dataout<=18'h04292;
					11'h0720: dataout<=18'h1f008;
					11'h0721: dataout<=18'h07ed9;
					11'h0722: dataout<=18'h1fbfd;
					11'h0723: dataout<=18'h03fec;
					11'h0724: dataout<=18'h1f154;
					11'h0725: dataout<=18'h079ab;
					11'h0726: dataout<=18'h1fc50;
					11'h0727: dataout<=18'h03d46;
					11'h0728: dataout<=18'h1f292;
					11'h0729: dataout<=18'h0747a;
					11'h072a: dataout<=18'h1fca0;
					11'h072b: dataout<=18'h03a9f;
					11'h072c: dataout<=18'h1f3c2;
					11'h072d: dataout<=18'h06f45;
					11'h072e: dataout<=18'h1fced;
					11'h072f: dataout<=18'h037f8;
					11'h0730: dataout<=18'h1f4e4;
					11'h0731: dataout<=18'h06a0e;
					11'h0732: dataout<=18'h1fd36;
					11'h0733: dataout<=18'h03551;
					11'h0734: dataout<=18'h1f5f8;
					11'h0735: dataout<=18'h064d3;
					11'h0736: dataout<=18'h1fd7b;
					11'h0737: dataout<=18'h032a9;
					11'h0738: dataout<=18'h1f6fe;
					11'h0739: dataout<=18'h05f95;
					11'h073a: dataout<=18'h1fdbd;
					11'h073b: dataout<=18'h03001;
					11'h073c: dataout<=18'h1f7f6;
					11'h073d: dataout<=18'h05a55;
					11'h073e: dataout<=18'h1fdfb;
					11'h073f: dataout<=18'h02d58;
					11'h0740: dataout<=18'h1f8e0;
					11'h0741: dataout<=18'h05513;
					11'h0742: dataout<=18'h1fe36;
					11'h0743: dataout<=18'h02aaf;
					11'h0744: dataout<=18'h1f9bc;
					11'h0745: dataout<=18'h04fce;
					11'h0746: dataout<=18'h1fe6d;
					11'h0747: dataout<=18'h02806;
					11'h0748: dataout<=18'h1fa8a;
					11'h0749: dataout<=18'h04a87;
					11'h074a: dataout<=18'h1fea1;
					11'h074b: dataout<=18'h0255d;
					11'h074c: dataout<=18'h1fb4a;
					11'h074d: dataout<=18'h0453d;
					11'h074e: dataout<=18'h1fed1;
					11'h074f: dataout<=18'h022b3;
					11'h0750: dataout<=18'h1fbfc;
					11'h0751: dataout<=18'h03ff2;
					11'h0752: dataout<=18'h1fefe;
					11'h0753: dataout<=18'h02009;
					11'h0754: dataout<=18'h1fca0;
					11'h0755: dataout<=18'h03aa5;
					11'h0756: dataout<=18'h1ff27;
					11'h0757: dataout<=18'h01d5f;
					11'h0758: dataout<=18'h1fd35;
					11'h0759: dataout<=18'h03556;
					11'h075a: dataout<=18'h1ff4c;
					11'h075b: dataout<=18'h01ab4;
					11'h075c: dataout<=18'h1fdbd;
					11'h075d: dataout<=18'h03006;
					11'h075e: dataout<=18'h1ff6e;
					11'h075f: dataout<=18'h0180a;
					11'h0760: dataout<=18'h1fe36;
					11'h0761: dataout<=18'h02ab5;
					11'h0762: dataout<=18'h1ff8c;
					11'h0763: dataout<=18'h0155f;
					11'h0764: dataout<=18'h1fea1;
					11'h0765: dataout<=18'h02562;
					11'h0766: dataout<=18'h1ffa7;
					11'h0767: dataout<=18'h012b4;
					11'h0768: dataout<=18'h1fefd;
					11'h0769: dataout<=18'h0200f;
					11'h076a: dataout<=18'h1ffbe;
					11'h076b: dataout<=18'h01009;
					11'h076c: dataout<=18'h1ff4c;
					11'h076d: dataout<=18'h01aba;
					11'h076e: dataout<=18'h1ffd2;
					11'h076f: dataout<=18'h00d5e;
					11'h0770: dataout<=18'h1ff8c;
					11'h0771: dataout<=18'h01565;
					11'h0772: dataout<=18'h1ffe2;
					11'h0773: dataout<=18'h00ab3;
					11'h0774: dataout<=18'h1ffbe;
					11'h0775: dataout<=18'h0100f;
					11'h0776: dataout<=18'h1ffee;
					11'h0777: dataout<=18'h00807;
					11'h0778: dataout<=18'h1ffe2;
					11'h0779: dataout<=18'h00ab8;
					11'h077a: dataout<=18'h1fff7;
					11'h077b: dataout<=18'h0055c;
					11'h077c: dataout<=18'h1ffe2;
					11'h077d: dataout<=18'h00ab8;
					11'h077e: dataout<=18'h1fff7;
					11'h077f: dataout<=18'h0055c;
					11'h0780: dataout<=18'h00000;
					11'h0781: dataout<=18'h00000;
					11'h0782: dataout<=18'h00000;
					11'h0783: dataout<=18'h00000;
					11'h0784: dataout<=18'h00000;
					11'h0785: dataout<=18'h00000;
					11'h0786: dataout<=18'h00000;
					11'h0787: dataout<=18'h00000;
					11'h0788: dataout<=18'h00000;
					11'h0789: dataout<=18'h00000;
					11'h078a: dataout<=18'h00000;
					11'h078b: dataout<=18'h00000;
					11'h078c: dataout<=18'h00000;
					11'h078d: dataout<=18'h00000;
					11'h078e: dataout<=18'h00000;
					11'h078f: dataout<=18'h00000;
					11'h0790: dataout<=18'h00000;
					11'h0791: dataout<=18'h00000;
					11'h0792: dataout<=18'h00000;
					11'h0793: dataout<=18'h00000;
					11'h0794: dataout<=18'h00000;
					11'h0795: dataout<=18'h00000;
					11'h0796: dataout<=18'h00000;
					11'h0797: dataout<=18'h00000;
					11'h0798: dataout<=18'h00000;
					11'h0799: dataout<=18'h00000;
					11'h079a: dataout<=18'h00000;
					11'h079b: dataout<=18'h00000;
					11'h079c: dataout<=18'h00000;
					11'h079d: dataout<=18'h00000;
					11'h079e: dataout<=18'h00000;
					11'h079f: dataout<=18'h00000;
					11'h07a0: dataout<=18'h00000;
					11'h07a1: dataout<=18'h00000;
					11'h07a2: dataout<=18'h00000;
					11'h07a3: dataout<=18'h00000;
					11'h07a4: dataout<=18'h00000;
					11'h07a5: dataout<=18'h00000;
					11'h07a6: dataout<=18'h00000;
					11'h07a7: dataout<=18'h00000;
					11'h07a8: dataout<=18'h00000;
					11'h07a9: dataout<=18'h00000;
					11'h07aa: dataout<=18'h00000;
					11'h07ab: dataout<=18'h00000;
					11'h07ac: dataout<=18'h00000;
					11'h07ad: dataout<=18'h00000;
					11'h07ae: dataout<=18'h00000;
					11'h07af: dataout<=18'h00000;
					11'h07b0: dataout<=18'h00000;
					11'h07b1: dataout<=18'h00000;
					11'h07b2: dataout<=18'h00000;
					11'h07b3: dataout<=18'h00000;
					11'h07b4: dataout<=18'h00000;
					11'h07b5: dataout<=18'h00000;
					11'h07b6: dataout<=18'h00000;
					11'h07b7: dataout<=18'h00000;
					11'h07b8: dataout<=18'h00000;
					11'h07b9: dataout<=18'h00000;
					11'h07ba: dataout<=18'h00000;
					11'h07bb: dataout<=18'h00000;
					11'h07bc: dataout<=18'h00000;
					11'h07bd: dataout<=18'h00000;
					11'h07be: dataout<=18'h00000;
					11'h07bf: dataout<=18'h00000;
					11'h07c0: dataout<=18'h00000;
					11'h07c1: dataout<=18'h00000;
					11'h07c2: dataout<=18'h00000;
					11'h07c3: dataout<=18'h00000;
					11'h07c4: dataout<=18'h00000;
					11'h07c5: dataout<=18'h00000;
					11'h07c6: dataout<=18'h00000;
					11'h07c7: dataout<=18'h00000;
					11'h07c8: dataout<=18'h00000;
					11'h07c9: dataout<=18'h00000;
					11'h07ca: dataout<=18'h00000;
					11'h07cb: dataout<=18'h00000;
					11'h07cc: dataout<=18'h00000;
					11'h07cd: dataout<=18'h00000;
					11'h07ce: dataout<=18'h00000;
					11'h07cf: dataout<=18'h00000;
					11'h07d0: dataout<=18'h00000;
					11'h07d1: dataout<=18'h00000;
					11'h07d2: dataout<=18'h00000;
					11'h07d3: dataout<=18'h00000;
					11'h07d4: dataout<=18'h00000;
					11'h07d5: dataout<=18'h00000;
					11'h07d6: dataout<=18'h00000;
					11'h07d7: dataout<=18'h00000;
					11'h07d8: dataout<=18'h00000;
					11'h07d9: dataout<=18'h00000;
					11'h07da: dataout<=18'h00000;
					11'h07db: dataout<=18'h00000;
					11'h07dc: dataout<=18'h00000;
					11'h07dd: dataout<=18'h00000;
					11'h07de: dataout<=18'h00000;
					11'h07df: dataout<=18'h00000;
					11'h07e0: dataout<=18'h00000;
					11'h07e1: dataout<=18'h00000;
					11'h07e2: dataout<=18'h00000;
					11'h07e3: dataout<=18'h00000;
					11'h07e4: dataout<=18'h00000;
					11'h07e5: dataout<=18'h00000;
					11'h07e6: dataout<=18'h00000;
					11'h07e7: dataout<=18'h00000;
					11'h07e8: dataout<=18'h00000;
					11'h07e9: dataout<=18'h00000;
					11'h07ea: dataout<=18'h00000;
					11'h07eb: dataout<=18'h00000;
					11'h07ec: dataout<=18'h00000;
					11'h07ed: dataout<=18'h00000;
					11'h07ee: dataout<=18'h00000;
					11'h07ef: dataout<=18'h00000;
					11'h07f0: dataout<=18'h00000;
					11'h07f1: dataout<=18'h00000;
					11'h07f2: dataout<=18'h00000;
					11'h07f3: dataout<=18'h00000;
					11'h07f4: dataout<=18'h00000;
					11'h07f5: dataout<=18'h00000;
					11'h07f6: dataout<=18'h00000;
					11'h07f7: dataout<=18'h00000;
					11'h07f8: dataout<=18'h00000;
					11'h07f9: dataout<=18'h00000;
					11'h07fa: dataout<=18'h00000;
					11'h07fb: dataout<=18'h00000;
					11'h07fc: dataout<=18'h00000;
					11'h07fd: dataout<=18'h00000;
					11'h07fe: dataout<=18'h00000;
					11'h07ff: dataout<=18'h00000;
				endcase
			end
		end
	end
endmodule

