module fctheta_rom (clock,ce,oce,reset,addr,dataout);
	input clock,ce,oce,reset;
	input [9:0] addr;
	output [35:0] dataout;
	reg [35:0] dataout;
	always @(posedge clock or posedge reset) begin
		if(reset) begin
			dataout <= 0;
		end else begin
			if (ce & oce) begin
				case (addr)
					10'd0000: dataout<=36'd27373258233;
					10'd0001: dataout<=36'd27316231610;
					10'd0002: dataout<=36'd27259204987;
					10'd0003: dataout<=36'd27202178364;
					10'd0004: dataout<=36'd27145151741;
					10'd0005: dataout<=36'd27088125118;
					10'd0006: dataout<=36'd27031098495;
					10'd0007: dataout<=36'd26974071872;
					10'd0008: dataout<=36'd26917045249;
					10'd0009: dataout<=36'd26860018626;
					10'd0010: dataout<=36'd26802992003;
					10'd0011: dataout<=36'd26745965380;
					10'd0012: dataout<=36'd26688938757;
					10'd0013: dataout<=36'd26631912134;
					10'd0014: dataout<=36'd26574885511;
					10'd0015: dataout<=36'd26517858888;
					10'd0016: dataout<=36'd26460832265;
					10'd0017: dataout<=36'd26403805642;
					10'd0018: dataout<=36'd26346779020;
					10'd0019: dataout<=36'd26289752397;
					10'd0020: dataout<=36'd26232725774;
					10'd0021: dataout<=36'd26175699151;
					10'd0022: dataout<=36'd26118672528;
					10'd0023: dataout<=36'd26061645905;
					10'd0024: dataout<=36'd26004619282;
					10'd0025: dataout<=36'd25947592659;
					10'd0026: dataout<=36'd25890566036;
					10'd0027: dataout<=36'd25833539413;
					10'd0028: dataout<=36'd25776512790;
					10'd0029: dataout<=36'd25719486167;
					10'd0030: dataout<=36'd25662459544;
					10'd0031: dataout<=36'd25605432921;
					10'd0032: dataout<=36'd25548406298;
					10'd0033: dataout<=36'd25491379675;
					10'd0034: dataout<=36'd25434353052;
					10'd0035: dataout<=36'd25377326429;
					10'd0036: dataout<=36'd25320299806;
					10'd0037: dataout<=36'd25263273183;
					10'd0038: dataout<=36'd25206246560;
					10'd0039: dataout<=36'd25149219937;
					10'd0040: dataout<=36'd25092193315;
					10'd0041: dataout<=36'd25035166692;
					10'd0042: dataout<=36'd24978140069;
					10'd0043: dataout<=36'd24921113446;
					10'd0044: dataout<=36'd24864086823;
					10'd0045: dataout<=36'd24807060200;
					10'd0046: dataout<=36'd24750033577;
					10'd0047: dataout<=36'd24693006954;
					10'd0048: dataout<=36'd24635980331;
					10'd0049: dataout<=36'd24578953708;
					10'd0050: dataout<=36'd24521927085;
					10'd0051: dataout<=36'd24464900462;
					10'd0052: dataout<=36'd24407873839;
					10'd0053: dataout<=36'd24350847216;
					10'd0054: dataout<=36'd24293820593;
					10'd0055: dataout<=36'd24236793970;
					10'd0056: dataout<=36'd24179767347;
					10'd0057: dataout<=36'd24122740724;
					10'd0058: dataout<=36'd24065714101;
					10'd0059: dataout<=36'd24008687478;
					10'd0060: dataout<=36'd23951660855;
					10'd0061: dataout<=36'd23894634232;
					10'd0062: dataout<=36'd23837607610;
					10'd0063: dataout<=36'd23780580987;
					10'd0064: dataout<=36'd23723554364;
					10'd0065: dataout<=36'd23666527741;
					10'd0066: dataout<=36'd23609501118;
					10'd0067: dataout<=36'd23552474495;
					10'd0068: dataout<=36'd23495447872;
					10'd0069: dataout<=36'd23438421249;
					10'd0070: dataout<=36'd23381394626;
					10'd0071: dataout<=36'd23324368003;
					10'd0072: dataout<=36'd23267341380;
					10'd0073: dataout<=36'd23210314757;
					10'd0074: dataout<=36'd23153288134;
					10'd0075: dataout<=36'd23096261511;
					10'd0076: dataout<=36'd23039234888;
					10'd0077: dataout<=36'd22982208265;
					10'd0078: dataout<=36'd22925181642;
					10'd0079: dataout<=36'd22868155019;
					10'd0080: dataout<=36'd22811128396;
					10'd0081: dataout<=36'd22754101773;
					10'd0082: dataout<=36'd22697075150;
					10'd0083: dataout<=36'd22640048528;
					10'd0084: dataout<=36'd22583021905;
					10'd0085: dataout<=36'd22525995282;
					10'd0086: dataout<=36'd22468968659;
					10'd0087: dataout<=36'd22411942036;
					10'd0088: dataout<=36'd22354915413;
					10'd0089: dataout<=36'd22297888790;
					10'd0090: dataout<=36'd22240862167;
					10'd0091: dataout<=36'd22183835544;
					10'd0092: dataout<=36'd22126808921;
					10'd0093: dataout<=36'd22069782298;
					10'd0094: dataout<=36'd22012755675;
					10'd0095: dataout<=36'd21955729052;
					10'd0096: dataout<=36'd21898702429;
					10'd0097: dataout<=36'd21841675806;
					10'd0098: dataout<=36'd21784649183;
					10'd0099: dataout<=36'd21727622560;
					10'd0100: dataout<=36'd21670595937;
					10'd0101: dataout<=36'd21613569314;
					10'd0102: dataout<=36'd21556542691;
					10'd0103: dataout<=36'd21499516068;
					10'd0104: dataout<=36'd21442489445;
					10'd0105: dataout<=36'd21385462823;
					10'd0106: dataout<=36'd21328436200;
					10'd0107: dataout<=36'd21271409577;
					10'd0108: dataout<=36'd21214382954;
					10'd0109: dataout<=36'd21157356331;
					10'd0110: dataout<=36'd21100329708;
					10'd0111: dataout<=36'd21043303085;
					10'd0112: dataout<=36'd20986276462;
					10'd0113: dataout<=36'd20929249839;
					10'd0114: dataout<=36'd20872223216;
					10'd0115: dataout<=36'd20815196593;
					10'd0116: dataout<=36'd20758169970;
					10'd0117: dataout<=36'd20701143347;
					10'd0118: dataout<=36'd20644116724;
					10'd0119: dataout<=36'd20587090101;
					10'd0120: dataout<=36'd20530063478;
					10'd0121: dataout<=36'd20473036855;
					10'd0122: dataout<=36'd20416010232;
					10'd0123: dataout<=36'd20358983609;
					10'd0124: dataout<=36'd20301956986;
					10'd0125: dataout<=36'd20244930363;
					10'd0126: dataout<=36'd20187903740;
					10'd0127: dataout<=36'd20130877118;
					10'd0128: dataout<=36'd20073850495;
					10'd0129: dataout<=36'd20016823872;
					10'd0130: dataout<=36'd19959797249;
					10'd0131: dataout<=36'd19902770626;
					10'd0132: dataout<=36'd19845744003;
					10'd0133: dataout<=36'd19788717380;
					10'd0134: dataout<=36'd19731690757;
					10'd0135: dataout<=36'd19674664134;
					10'd0136: dataout<=36'd19617637511;
					10'd0137: dataout<=36'd19560610888;
					10'd0138: dataout<=36'd19503584265;
					10'd0139: dataout<=36'd19446557642;
					10'd0140: dataout<=36'd19389531019;
					10'd0141: dataout<=36'd19332504396;
					10'd0142: dataout<=36'd19275477773;
					10'd0143: dataout<=36'd19218451150;
					10'd0144: dataout<=36'd19161424527;
					10'd0145: dataout<=36'd19104397904;
					10'd0146: dataout<=36'd19047371281;
					10'd0147: dataout<=36'd18990344658;
					10'd0148: dataout<=36'd18933318036;
					10'd0149: dataout<=36'd18876291413;
					10'd0150: dataout<=36'd18819264790;
					10'd0151: dataout<=36'd18762238167;
					10'd0152: dataout<=36'd18705211544;
					10'd0153: dataout<=36'd18648184921;
					10'd0154: dataout<=36'd18591158298;
					10'd0155: dataout<=36'd18534131675;
					10'd0156: dataout<=36'd18477105052;
					10'd0157: dataout<=36'd18420078429;
					10'd0158: dataout<=36'd18363051806;
					10'd0159: dataout<=36'd18306025183;
					10'd0160: dataout<=36'd18248998560;
					10'd0161: dataout<=36'd18191971937;
					10'd0162: dataout<=36'd18134945314;
					10'd0163: dataout<=36'd18077918691;
					10'd0164: dataout<=36'd18020892068;
					10'd0165: dataout<=36'd17963865445;
					10'd0166: dataout<=36'd17906838822;
					10'd0167: dataout<=36'd17849812199;
					10'd0168: dataout<=36'd17792785576;
					10'd0169: dataout<=36'd17735758953;
					10'd0170: dataout<=36'd17678732331;
					10'd0171: dataout<=36'd17621705708;
					10'd0172: dataout<=36'd17564679085;
					10'd0173: dataout<=36'd17507652462;
					10'd0174: dataout<=36'd17450625839;
					10'd0175: dataout<=36'd17393599216;
					10'd0176: dataout<=36'd17336572593;
					10'd0177: dataout<=36'd17279545970;
					10'd0178: dataout<=36'd17222519347;
					10'd0179: dataout<=36'd17165492724;
					10'd0180: dataout<=36'd17108466101;
					10'd0181: dataout<=36'd17051439478;
					10'd0182: dataout<=36'd16994412855;
					10'd0183: dataout<=36'd16937386232;
					10'd0184: dataout<=36'd16880359609;
					10'd0185: dataout<=36'd16823332986;
					10'd0186: dataout<=36'd16766306363;
					10'd0187: dataout<=36'd16709279740;
					10'd0188: dataout<=36'd16652253117;
					10'd0189: dataout<=36'd16595226494;
					10'd0190: dataout<=36'd16538199871;
					10'd0191: dataout<=36'd16481173248;
					10'd0192: dataout<=36'd16424146626;
					10'd0193: dataout<=36'd16367120003;
					10'd0194: dataout<=36'd16310093380;
					10'd0195: dataout<=36'd16253066757;
					10'd0196: dataout<=36'd16196040134;
					10'd0197: dataout<=36'd16139013511;
					10'd0198: dataout<=36'd16081986888;
					10'd0199: dataout<=36'd16024960265;
					10'd0200: dataout<=36'd15967933642;
					10'd0201: dataout<=36'd15910907019;
					10'd0202: dataout<=36'd15853880396;
					10'd0203: dataout<=36'd15796853773;
					10'd0204: dataout<=36'd15739827150;
					10'd0205: dataout<=36'd15682800527;
					10'd0206: dataout<=36'd15625773904;
					10'd0207: dataout<=36'd15568747281;
					10'd0208: dataout<=36'd15511720658;
					10'd0209: dataout<=36'd15454694035;
					10'd0210: dataout<=36'd15397667412;
					10'd0211: dataout<=36'd15340640789;
					10'd0212: dataout<=36'd15283614166;
					10'd0213: dataout<=36'd15226587544;
					10'd0214: dataout<=36'd15169560921;
					10'd0215: dataout<=36'd15112534298;
					10'd0216: dataout<=36'd15055507675;
					10'd0217: dataout<=36'd14998481052;
					10'd0218: dataout<=36'd14941454429;
					10'd0219: dataout<=36'd14884427806;
					10'd0220: dataout<=36'd14827401183;
					10'd0221: dataout<=36'd14770374560;
					10'd0222: dataout<=36'd14713347937;
					10'd0223: dataout<=36'd14656321314;
					10'd0224: dataout<=36'd14599294691;
					10'd0225: dataout<=36'd14542268068;
					10'd0226: dataout<=36'd14485241445;
					10'd0227: dataout<=36'd14428214822;
					10'd0228: dataout<=36'd14371188199;
					10'd0229: dataout<=36'd14314161576;
					10'd0230: dataout<=36'd14257134953;
					10'd0231: dataout<=36'd14200108330;
					10'd0232: dataout<=36'd14143081707;
					10'd0233: dataout<=36'd14086055084;
					10'd0234: dataout<=36'd14029028461;
					10'd0235: dataout<=36'd13972001839;
					10'd0236: dataout<=36'd13914975216;
					10'd0237: dataout<=36'd13857948593;
					10'd0238: dataout<=36'd13800921970;
					10'd0239: dataout<=36'd13743895347;
					10'd0240: dataout<=36'd13686868724;
					10'd0241: dataout<=36'd13629842101;
					10'd0242: dataout<=36'd13572815478;
					10'd0243: dataout<=36'd13515788855;
					10'd0244: dataout<=36'd13458762232;
					10'd0245: dataout<=36'd13401735609;
					10'd0246: dataout<=36'd13344708986;
					10'd0247: dataout<=36'd13287682363;
					10'd0248: dataout<=36'd13230655740;
					10'd0249: dataout<=36'd13173629117;
					10'd0250: dataout<=36'd13116602494;
					10'd0251: dataout<=36'd13059575871;
					10'd0252: dataout<=36'd13002549248;
					10'd0253: dataout<=36'd12945522625;
					10'd0254: dataout<=36'd12888496002;
					10'd0255: dataout<=36'd12831469379;
					10'd0256: dataout<=36'd12774442756;
					10'd0257: dataout<=36'd12717416134;
					10'd0258: dataout<=36'd12660389511;
					10'd0259: dataout<=36'd12603362888;
					10'd0260: dataout<=36'd12546336265;
					10'd0261: dataout<=36'd12489309642;
					10'd0262: dataout<=36'd12432283019;
					10'd0263: dataout<=36'd12375256396;
					10'd0264: dataout<=36'd12318229773;
					10'd0265: dataout<=36'd12261203150;
					10'd0266: dataout<=36'd12204176527;
					10'd0267: dataout<=36'd12147149904;
					10'd0268: dataout<=36'd12090123281;
					10'd0269: dataout<=36'd12033096658;
					10'd0270: dataout<=36'd11976070035;
					10'd0271: dataout<=36'd11919043412;
					10'd0272: dataout<=36'd11862016789;
					10'd0273: dataout<=36'd11804990166;
					10'd0274: dataout<=36'd11747963543;
					10'd0275: dataout<=36'd11690936920;
					10'd0276: dataout<=36'd11633910297;
					10'd0277: dataout<=36'd11576883674;
					10'd0278: dataout<=36'd11519857051;
					10'd0279: dataout<=36'd11462830429;
					10'd0280: dataout<=36'd11405803806;
					10'd0281: dataout<=36'd11348777183;
					10'd0282: dataout<=36'd11291750560;
					10'd0283: dataout<=36'd11234723937;
					10'd0284: dataout<=36'd11177697314;
					10'd0285: dataout<=36'd11120670691;
					10'd0286: dataout<=36'd11063644068;
					10'd0287: dataout<=36'd11006617445;
					10'd0288: dataout<=36'd10949590822;
					10'd0289: dataout<=36'd10892564199;
					10'd0290: dataout<=36'd10835537576;
					10'd0291: dataout<=36'd10778510953;
					10'd0292: dataout<=36'd10721484330;
					10'd0293: dataout<=36'd10664457707;
					10'd0294: dataout<=36'd10607431084;
					10'd0295: dataout<=36'd10550404461;
					10'd0296: dataout<=36'd10493377838;
					10'd0297: dataout<=36'd10436351215;
					10'd0298: dataout<=36'd10379324592;
					10'd0299: dataout<=36'd10322297969;
					10'd0300: dataout<=36'd10265271347;
					10'd0301: dataout<=36'd10208244724;
					10'd0302: dataout<=36'd10151218101;
					10'd0303: dataout<=36'd10094191478;
					10'd0304: dataout<=36'd10037164855;
					10'd0305: dataout<=36'd9980138232;
					10'd0306: dataout<=36'd9923111609;
					10'd0307: dataout<=36'd9866084986;
					10'd0308: dataout<=36'd9809058363;
					10'd0309: dataout<=36'd9752031740;
					10'd0310: dataout<=36'd9695005117;
					10'd0311: dataout<=36'd9637978494;
					10'd0312: dataout<=36'd9580951871;
					10'd0313: dataout<=36'd9523925248;
					10'd0314: dataout<=36'd9466898625;
					10'd0315: dataout<=36'd9409872002;
					10'd0316: dataout<=36'd9352845379;
					10'd0317: dataout<=36'd9295818756;
					10'd0318: dataout<=36'd9238792133;
					10'd0319: dataout<=36'd9181765510;
					10'd0320: dataout<=36'd9124738887;
					10'd0321: dataout<=36'd9067712264;
					10'd0322: dataout<=36'd9010685642;
					10'd0323: dataout<=36'd8953659019;
					10'd0324: dataout<=36'd8896632396;
					10'd0325: dataout<=36'd8839605773;
					10'd0326: dataout<=36'd8782579150;
					10'd0327: dataout<=36'd8725552527;
					10'd0328: dataout<=36'd8668525904;
					10'd0329: dataout<=36'd8611499281;
					10'd0330: dataout<=36'd8554472658;
					10'd0331: dataout<=36'd8497446035;
					10'd0332: dataout<=36'd8440419412;
					10'd0333: dataout<=36'd8383392789;
					10'd0334: dataout<=36'd8326366166;
					10'd0335: dataout<=36'd8269339543;
					10'd0336: dataout<=36'd8212312920;
					10'd0337: dataout<=36'd8155286297;
					10'd0338: dataout<=36'd8098259674;
					10'd0339: dataout<=36'd8041233051;
					10'd0340: dataout<=36'd7984206428;
					10'd0341: dataout<=36'd7927179805;
					10'd0342: dataout<=36'd7870153182;
					10'd0343: dataout<=36'd7813126559;
					10'd0344: dataout<=36'd7756099937;
					10'd0345: dataout<=36'd7699073314;
					10'd0346: dataout<=36'd7642046691;
					10'd0347: dataout<=36'd7585020068;
					10'd0348: dataout<=36'd7527993445;
					10'd0349: dataout<=36'd7470966822;
					10'd0350: dataout<=36'd7413940199;
					10'd0351: dataout<=36'd7356913576;
					10'd0352: dataout<=36'd7299886953;
					10'd0353: dataout<=36'd7242860330;
					10'd0354: dataout<=36'd7185833707;
					10'd0355: dataout<=36'd7128807084;
					10'd0356: dataout<=36'd7071780461;
					10'd0357: dataout<=36'd7014753838;
					10'd0358: dataout<=36'd6957727215;
					10'd0359: dataout<=36'd6900700592;
					10'd0360: dataout<=36'd6843673969;
					10'd0361: dataout<=36'd6786647346;
					10'd0362: dataout<=36'd6729620723;
					10'd0363: dataout<=36'd6672594100;
					10'd0364: dataout<=36'd6615567477;
					10'd0365: dataout<=36'd6558540855;
					10'd0366: dataout<=36'd6501514232;
					10'd0367: dataout<=36'd6444487609;
					10'd0368: dataout<=36'd6387460986;
					10'd0369: dataout<=36'd6330434363;
					10'd0370: dataout<=36'd6273407740;
					10'd0371: dataout<=36'd6216381117;
					10'd0372: dataout<=36'd6159354494;
					10'd0373: dataout<=36'd6102327871;
					10'd0374: dataout<=36'd6045301248;
					10'd0375: dataout<=36'd5988274625;
					10'd0376: dataout<=36'd5931248002;
					10'd0377: dataout<=36'd5874221379;
					10'd0378: dataout<=36'd5817194756;
					10'd0379: dataout<=36'd5760168133;
					10'd0380: dataout<=36'd5703141510;
					10'd0381: dataout<=36'd5646114887;
					10'd0382: dataout<=36'd5589088264;
					10'd0383: dataout<=36'd5532061641;
					10'd0384: dataout<=36'd5475035018;
					10'd0385: dataout<=36'd5418008395;
					10'd0386: dataout<=36'd5360981772;
					10'd0387: dataout<=36'd5303955150;
					10'd0388: dataout<=36'd5246928527;
					10'd0389: dataout<=36'd5189901904;
					10'd0390: dataout<=36'd5132875281;
					10'd0391: dataout<=36'd5075848658;
					10'd0392: dataout<=36'd5018822035;
					10'd0393: dataout<=36'd4961795412;
					10'd0394: dataout<=36'd4904768789;
					10'd0395: dataout<=36'd4847742166;
					10'd0396: dataout<=36'd4790715543;
					10'd0397: dataout<=36'd4733688920;
					10'd0398: dataout<=36'd4676662297;
					10'd0399: dataout<=36'd4619635674;
					10'd0400: dataout<=36'd4562609051;
					10'd0401: dataout<=36'd4505582428;
					10'd0402: dataout<=36'd4448555805;
					10'd0403: dataout<=36'd4391529182;
					10'd0404: dataout<=36'd4334502559;
					10'd0405: dataout<=36'd4277475936;
					10'd0406: dataout<=36'd4220449313;
					10'd0407: dataout<=36'd4163422690;
					10'd0408: dataout<=36'd4106396067;
					10'd0409: dataout<=36'd4049369445;
					10'd0410: dataout<=36'd3992342822;
					10'd0411: dataout<=36'd3935316199;
					10'd0412: dataout<=36'd3878289576;
					10'd0413: dataout<=36'd3821262953;
					10'd0414: dataout<=36'd3764236330;
					10'd0415: dataout<=36'd3707209707;
					10'd0416: dataout<=36'd3650183084;
					10'd0417: dataout<=36'd3593156461;
					10'd0418: dataout<=36'd3536129838;
					10'd0419: dataout<=36'd3479103215;
					10'd0420: dataout<=36'd3422076592;
					10'd0421: dataout<=36'd3365049969;
					10'd0422: dataout<=36'd3308023346;
					10'd0423: dataout<=36'd3250996723;
					10'd0424: dataout<=36'd3193970100;
					10'd0425: dataout<=36'd3136943477;
					10'd0426: dataout<=36'd3079916854;
					10'd0427: dataout<=36'd3022890231;
					10'd0428: dataout<=36'd2965863608;
					10'd0429: dataout<=36'd2908836985;
					10'd0430: dataout<=36'd2851810363;
					10'd0431: dataout<=36'd2794783740;
					10'd0432: dataout<=36'd2737757117;
					10'd0433: dataout<=36'd2680730494;
					10'd0434: dataout<=36'd2623703871;
					10'd0435: dataout<=36'd2566677248;
					10'd0436: dataout<=36'd2509650625;
					10'd0437: dataout<=36'd2452624002;
					10'd0438: dataout<=36'd2395597379;
					10'd0439: dataout<=36'd2338570756;
					10'd0440: dataout<=36'd2281544133;
					10'd0441: dataout<=36'd2224517510;
					10'd0442: dataout<=36'd2167490887;
					10'd0443: dataout<=36'd2110464264;
					10'd0444: dataout<=36'd2053437641;
					10'd0445: dataout<=36'd1996411018;
					10'd0446: dataout<=36'd1939384395;
					10'd0447: dataout<=36'd1882357772;
					10'd0448: dataout<=36'd1825331149;
					10'd0449: dataout<=36'd1768304526;
					10'd0450: dataout<=36'd1711277903;
					10'd0451: dataout<=36'd1654251280;
					10'd0452: dataout<=36'd1597224658;
					10'd0453: dataout<=36'd1540198035;
					10'd0454: dataout<=36'd1483171412;
					10'd0455: dataout<=36'd1426144789;
					10'd0456: dataout<=36'd1369118166;
					10'd0457: dataout<=36'd1312091543;
					10'd0458: dataout<=36'd1255064920;
					10'd0459: dataout<=36'd1198038297;
					10'd0460: dataout<=36'd1141011674;
					10'd0461: dataout<=36'd1083985051;
					10'd0462: dataout<=36'd1026958428;
					10'd0463: dataout<=36'd969931805;
					10'd0464: dataout<=36'd912905182;
					10'd0465: dataout<=36'd855878559;
					10'd0466: dataout<=36'd798851936;
					10'd0467: dataout<=36'd741825313;
					10'd0468: dataout<=36'd684798690;
					10'd0469: dataout<=36'd627772067;
					10'd0470: dataout<=36'd570745444;
					10'd0471: dataout<=36'd513718821;
					10'd0472: dataout<=36'd456692198;
					10'd0473: dataout<=36'd399665575;
					10'd0474: dataout<=36'd342638953;
					10'd0475: dataout<=36'd285612330;
					10'd0476: dataout<=36'd228585707;
					10'd0477: dataout<=36'd171559084;
					10'd0478: dataout<=36'd114532461;
					10'd0479: dataout<=36'd114532461;
					10'd0480: dataout<=36'd00000000;
					10'd0481: dataout<=36'd00000000;
					10'd0482: dataout<=36'd00000000;
					10'd0483: dataout<=36'd00000000;
					10'd0484: dataout<=36'd00000000;
					10'd0485: dataout<=36'd00000000;
					10'd0486: dataout<=36'd00000000;
					10'd0487: dataout<=36'd00000000;
					10'd0488: dataout<=36'd00000000;
					10'd0489: dataout<=36'd00000000;
					10'd0490: dataout<=36'd00000000;
					10'd0491: dataout<=36'd00000000;
					10'd0492: dataout<=36'd00000000;
					10'd0493: dataout<=36'd00000000;
					10'd0494: dataout<=36'd00000000;
					10'd0495: dataout<=36'd00000000;
					10'd0496: dataout<=36'd00000000;
					10'd0497: dataout<=36'd00000000;
					10'd0498: dataout<=36'd00000000;
					10'd0499: dataout<=36'd00000000;
					10'd0500: dataout<=36'd00000000;
					10'd0501: dataout<=36'd00000000;
					10'd0502: dataout<=36'd00000000;
					10'd0503: dataout<=36'd00000000;
					10'd0504: dataout<=36'd00000000;
					10'd0505: dataout<=36'd00000000;
					10'd0506: dataout<=36'd00000000;
					10'd0507: dataout<=36'd00000000;
					10'd0508: dataout<=36'd00000000;
					10'd0509: dataout<=36'd00000000;
					10'd0510: dataout<=36'd00000000;
					10'd0511: dataout<=36'd00000000;
					10'd0512: dataout<=36'd00000000;
					10'd0513: dataout<=36'd00000000;
					10'd0514: dataout<=36'd00000000;
					10'd0515: dataout<=36'd00000000;
					10'd0516: dataout<=36'd00000000;
					10'd0517: dataout<=36'd00000000;
					10'd0518: dataout<=36'd00000000;
					10'd0519: dataout<=36'd00000000;
					10'd0520: dataout<=36'd00000000;
					10'd0521: dataout<=36'd00000000;
					10'd0522: dataout<=36'd00000000;
					10'd0523: dataout<=36'd00000000;
					10'd0524: dataout<=36'd00000000;
					10'd0525: dataout<=36'd00000000;
					10'd0526: dataout<=36'd00000000;
					10'd0527: dataout<=36'd00000000;
					10'd0528: dataout<=36'd00000000;
					10'd0529: dataout<=36'd00000000;
					10'd0530: dataout<=36'd00000000;
					10'd0531: dataout<=36'd00000000;
					10'd0532: dataout<=36'd00000000;
					10'd0533: dataout<=36'd00000000;
					10'd0534: dataout<=36'd00000000;
					10'd0535: dataout<=36'd00000000;
					10'd0536: dataout<=36'd00000000;
					10'd0537: dataout<=36'd00000000;
					10'd0538: dataout<=36'd00000000;
					10'd0539: dataout<=36'd00000000;
					10'd0540: dataout<=36'd00000000;
					10'd0541: dataout<=36'd00000000;
					10'd0542: dataout<=36'd00000000;
					10'd0543: dataout<=36'd00000000;
					10'd0544: dataout<=36'd00000000;
					10'd0545: dataout<=36'd00000000;
					10'd0546: dataout<=36'd00000000;
					10'd0547: dataout<=36'd00000000;
					10'd0548: dataout<=36'd00000000;
					10'd0549: dataout<=36'd00000000;
					10'd0550: dataout<=36'd00000000;
					10'd0551: dataout<=36'd00000000;
					10'd0552: dataout<=36'd00000000;
					10'd0553: dataout<=36'd00000000;
					10'd0554: dataout<=36'd00000000;
					10'd0555: dataout<=36'd00000000;
					10'd0556: dataout<=36'd00000000;
					10'd0557: dataout<=36'd00000000;
					10'd0558: dataout<=36'd00000000;
					10'd0559: dataout<=36'd00000000;
					10'd0560: dataout<=36'd00000000;
					10'd0561: dataout<=36'd00000000;
					10'd0562: dataout<=36'd00000000;
					10'd0563: dataout<=36'd00000000;
					10'd0564: dataout<=36'd00000000;
					10'd0565: dataout<=36'd00000000;
					10'd0566: dataout<=36'd00000000;
					10'd0567: dataout<=36'd00000000;
					10'd0568: dataout<=36'd00000000;
					10'd0569: dataout<=36'd00000000;
					10'd0570: dataout<=36'd00000000;
					10'd0571: dataout<=36'd00000000;
					10'd0572: dataout<=36'd00000000;
					10'd0573: dataout<=36'd00000000;
					10'd0574: dataout<=36'd00000000;
					10'd0575: dataout<=36'd00000000;
					10'd0576: dataout<=36'd00000000;
					10'd0577: dataout<=36'd00000000;
					10'd0578: dataout<=36'd00000000;
					10'd0579: dataout<=36'd00000000;
					10'd0580: dataout<=36'd00000000;
					10'd0581: dataout<=36'd00000000;
					10'd0582: dataout<=36'd00000000;
					10'd0583: dataout<=36'd00000000;
					10'd0584: dataout<=36'd00000000;
					10'd0585: dataout<=36'd00000000;
					10'd0586: dataout<=36'd00000000;
					10'd0587: dataout<=36'd00000000;
					10'd0588: dataout<=36'd00000000;
					10'd0589: dataout<=36'd00000000;
					10'd0590: dataout<=36'd00000000;
					10'd0591: dataout<=36'd00000000;
					10'd0592: dataout<=36'd00000000;
					10'd0593: dataout<=36'd00000000;
					10'd0594: dataout<=36'd00000000;
					10'd0595: dataout<=36'd00000000;
					10'd0596: dataout<=36'd00000000;
					10'd0597: dataout<=36'd00000000;
					10'd0598: dataout<=36'd00000000;
					10'd0599: dataout<=36'd00000000;
					10'd0600: dataout<=36'd00000000;
					10'd0601: dataout<=36'd00000000;
					10'd0602: dataout<=36'd00000000;
					10'd0603: dataout<=36'd00000000;
					10'd0604: dataout<=36'd00000000;
					10'd0605: dataout<=36'd00000000;
					10'd0606: dataout<=36'd00000000;
					10'd0607: dataout<=36'd00000000;
					10'd0608: dataout<=36'd00000000;
					10'd0609: dataout<=36'd00000000;
					10'd0610: dataout<=36'd00000000;
					10'd0611: dataout<=36'd00000000;
					10'd0612: dataout<=36'd00000000;
					10'd0613: dataout<=36'd00000000;
					10'd0614: dataout<=36'd00000000;
					10'd0615: dataout<=36'd00000000;
					10'd0616: dataout<=36'd00000000;
					10'd0617: dataout<=36'd00000000;
					10'd0618: dataout<=36'd00000000;
					10'd0619: dataout<=36'd00000000;
					10'd0620: dataout<=36'd00000000;
					10'd0621: dataout<=36'd00000000;
					10'd0622: dataout<=36'd00000000;
					10'd0623: dataout<=36'd00000000;
					10'd0624: dataout<=36'd00000000;
					10'd0625: dataout<=36'd00000000;
					10'd0626: dataout<=36'd00000000;
					10'd0627: dataout<=36'd00000000;
					10'd0628: dataout<=36'd00000000;
					10'd0629: dataout<=36'd00000000;
					10'd0630: dataout<=36'd00000000;
					10'd0631: dataout<=36'd00000000;
					10'd0632: dataout<=36'd00000000;
					10'd0633: dataout<=36'd00000000;
					10'd0634: dataout<=36'd00000000;
					10'd0635: dataout<=36'd00000000;
					10'd0636: dataout<=36'd00000000;
					10'd0637: dataout<=36'd00000000;
					10'd0638: dataout<=36'd00000000;
					10'd0639: dataout<=36'd00000000;
					10'd0640: dataout<=36'd00000000;
					10'd0641: dataout<=36'd00000000;
					10'd0642: dataout<=36'd00000000;
					10'd0643: dataout<=36'd00000000;
					10'd0644: dataout<=36'd00000000;
					10'd0645: dataout<=36'd00000000;
					10'd0646: dataout<=36'd00000000;
					10'd0647: dataout<=36'd00000000;
					10'd0648: dataout<=36'd00000000;
					10'd0649: dataout<=36'd00000000;
					10'd0650: dataout<=36'd00000000;
					10'd0651: dataout<=36'd00000000;
					10'd0652: dataout<=36'd00000000;
					10'd0653: dataout<=36'd00000000;
					10'd0654: dataout<=36'd00000000;
					10'd0655: dataout<=36'd00000000;
					10'd0656: dataout<=36'd00000000;
					10'd0657: dataout<=36'd00000000;
					10'd0658: dataout<=36'd00000000;
					10'd0659: dataout<=36'd00000000;
					10'd0660: dataout<=36'd00000000;
					10'd0661: dataout<=36'd00000000;
					10'd0662: dataout<=36'd00000000;
					10'd0663: dataout<=36'd00000000;
					10'd0664: dataout<=36'd00000000;
					10'd0665: dataout<=36'd00000000;
					10'd0666: dataout<=36'd00000000;
					10'd0667: dataout<=36'd00000000;
					10'd0668: dataout<=36'd00000000;
					10'd0669: dataout<=36'd00000000;
					10'd0670: dataout<=36'd00000000;
					10'd0671: dataout<=36'd00000000;
					10'd0672: dataout<=36'd00000000;
					10'd0673: dataout<=36'd00000000;
					10'd0674: dataout<=36'd00000000;
					10'd0675: dataout<=36'd00000000;
					10'd0676: dataout<=36'd00000000;
					10'd0677: dataout<=36'd00000000;
					10'd0678: dataout<=36'd00000000;
					10'd0679: dataout<=36'd00000000;
					10'd0680: dataout<=36'd00000000;
					10'd0681: dataout<=36'd00000000;
					10'd0682: dataout<=36'd00000000;
					10'd0683: dataout<=36'd00000000;
					10'd0684: dataout<=36'd00000000;
					10'd0685: dataout<=36'd00000000;
					10'd0686: dataout<=36'd00000000;
					10'd0687: dataout<=36'd00000000;
					10'd0688: dataout<=36'd00000000;
					10'd0689: dataout<=36'd00000000;
					10'd0690: dataout<=36'd00000000;
					10'd0691: dataout<=36'd00000000;
					10'd0692: dataout<=36'd00000000;
					10'd0693: dataout<=36'd00000000;
					10'd0694: dataout<=36'd00000000;
					10'd0695: dataout<=36'd00000000;
					10'd0696: dataout<=36'd00000000;
					10'd0697: dataout<=36'd00000000;
					10'd0698: dataout<=36'd00000000;
					10'd0699: dataout<=36'd00000000;
					10'd0700: dataout<=36'd00000000;
					10'd0701: dataout<=36'd00000000;
					10'd0702: dataout<=36'd00000000;
					10'd0703: dataout<=36'd00000000;
					10'd0704: dataout<=36'd00000000;
					10'd0705: dataout<=36'd00000000;
					10'd0706: dataout<=36'd00000000;
					10'd0707: dataout<=36'd00000000;
					10'd0708: dataout<=36'd00000000;
					10'd0709: dataout<=36'd00000000;
					10'd0710: dataout<=36'd00000000;
					10'd0711: dataout<=36'd00000000;
					10'd0712: dataout<=36'd00000000;
					10'd0713: dataout<=36'd00000000;
					10'd0714: dataout<=36'd00000000;
					10'd0715: dataout<=36'd00000000;
					10'd0716: dataout<=36'd00000000;
					10'd0717: dataout<=36'd00000000;
					10'd0718: dataout<=36'd00000000;
					10'd0719: dataout<=36'd00000000;
					10'd0720: dataout<=36'd00000000;
					10'd0721: dataout<=36'd00000000;
					10'd0722: dataout<=36'd00000000;
					10'd0723: dataout<=36'd00000000;
					10'd0724: dataout<=36'd00000000;
					10'd0725: dataout<=36'd00000000;
					10'd0726: dataout<=36'd00000000;
					10'd0727: dataout<=36'd00000000;
					10'd0728: dataout<=36'd00000000;
					10'd0729: dataout<=36'd00000000;
					10'd0730: dataout<=36'd00000000;
					10'd0731: dataout<=36'd00000000;
					10'd0732: dataout<=36'd00000000;
					10'd0733: dataout<=36'd00000000;
					10'd0734: dataout<=36'd00000000;
					10'd0735: dataout<=36'd00000000;
					10'd0736: dataout<=36'd00000000;
					10'd0737: dataout<=36'd00000000;
					10'd0738: dataout<=36'd00000000;
					10'd0739: dataout<=36'd00000000;
					10'd0740: dataout<=36'd00000000;
					10'd0741: dataout<=36'd00000000;
					10'd0742: dataout<=36'd00000000;
					10'd0743: dataout<=36'd00000000;
					10'd0744: dataout<=36'd00000000;
					10'd0745: dataout<=36'd00000000;
					10'd0746: dataout<=36'd00000000;
					10'd0747: dataout<=36'd00000000;
					10'd0748: dataout<=36'd00000000;
					10'd0749: dataout<=36'd00000000;
					10'd0750: dataout<=36'd00000000;
					10'd0751: dataout<=36'd00000000;
					10'd0752: dataout<=36'd00000000;
					10'd0753: dataout<=36'd00000000;
					10'd0754: dataout<=36'd00000000;
					10'd0755: dataout<=36'd00000000;
					10'd0756: dataout<=36'd00000000;
					10'd0757: dataout<=36'd00000000;
					10'd0758: dataout<=36'd00000000;
					10'd0759: dataout<=36'd00000000;
					10'd0760: dataout<=36'd00000000;
					10'd0761: dataout<=36'd00000000;
					10'd0762: dataout<=36'd00000000;
					10'd0763: dataout<=36'd00000000;
					10'd0764: dataout<=36'd00000000;
					10'd0765: dataout<=36'd00000000;
					10'd0766: dataout<=36'd00000000;
					10'd0767: dataout<=36'd00000000;
					10'd0768: dataout<=36'd00000000;
					10'd0769: dataout<=36'd00000000;
					10'd0770: dataout<=36'd00000000;
					10'd0771: dataout<=36'd00000000;
					10'd0772: dataout<=36'd00000000;
					10'd0773: dataout<=36'd00000000;
					10'd0774: dataout<=36'd00000000;
					10'd0775: dataout<=36'd00000000;
					10'd0776: dataout<=36'd00000000;
					10'd0777: dataout<=36'd00000000;
					10'd0778: dataout<=36'd00000000;
					10'd0779: dataout<=36'd00000000;
					10'd0780: dataout<=36'd00000000;
					10'd0781: dataout<=36'd00000000;
					10'd0782: dataout<=36'd00000000;
					10'd0783: dataout<=36'd00000000;
					10'd0784: dataout<=36'd00000000;
					10'd0785: dataout<=36'd00000000;
					10'd0786: dataout<=36'd00000000;
					10'd0787: dataout<=36'd00000000;
					10'd0788: dataout<=36'd00000000;
					10'd0789: dataout<=36'd00000000;
					10'd0790: dataout<=36'd00000000;
					10'd0791: dataout<=36'd00000000;
					10'd0792: dataout<=36'd00000000;
					10'd0793: dataout<=36'd00000000;
					10'd0794: dataout<=36'd00000000;
					10'd0795: dataout<=36'd00000000;
					10'd0796: dataout<=36'd00000000;
					10'd0797: dataout<=36'd00000000;
					10'd0798: dataout<=36'd00000000;
					10'd0799: dataout<=36'd00000000;
					10'd0800: dataout<=36'd00000000;
					10'd0801: dataout<=36'd00000000;
					10'd0802: dataout<=36'd00000000;
					10'd0803: dataout<=36'd00000000;
					10'd0804: dataout<=36'd00000000;
					10'd0805: dataout<=36'd00000000;
					10'd0806: dataout<=36'd00000000;
					10'd0807: dataout<=36'd00000000;
					10'd0808: dataout<=36'd00000000;
					10'd0809: dataout<=36'd00000000;
					10'd0810: dataout<=36'd00000000;
					10'd0811: dataout<=36'd00000000;
					10'd0812: dataout<=36'd00000000;
					10'd0813: dataout<=36'd00000000;
					10'd0814: dataout<=36'd00000000;
					10'd0815: dataout<=36'd00000000;
					10'd0816: dataout<=36'd00000000;
					10'd0817: dataout<=36'd00000000;
					10'd0818: dataout<=36'd00000000;
					10'd0819: dataout<=36'd00000000;
					10'd0820: dataout<=36'd00000000;
					10'd0821: dataout<=36'd00000000;
					10'd0822: dataout<=36'd00000000;
					10'd0823: dataout<=36'd00000000;
					10'd0824: dataout<=36'd00000000;
					10'd0825: dataout<=36'd00000000;
					10'd0826: dataout<=36'd00000000;
					10'd0827: dataout<=36'd00000000;
					10'd0828: dataout<=36'd00000000;
					10'd0829: dataout<=36'd00000000;
					10'd0830: dataout<=36'd00000000;
					10'd0831: dataout<=36'd00000000;
					10'd0832: dataout<=36'd00000000;
					10'd0833: dataout<=36'd00000000;
					10'd0834: dataout<=36'd00000000;
					10'd0835: dataout<=36'd00000000;
					10'd0836: dataout<=36'd00000000;
					10'd0837: dataout<=36'd00000000;
					10'd0838: dataout<=36'd00000000;
					10'd0839: dataout<=36'd00000000;
					10'd0840: dataout<=36'd00000000;
					10'd0841: dataout<=36'd00000000;
					10'd0842: dataout<=36'd00000000;
					10'd0843: dataout<=36'd00000000;
					10'd0844: dataout<=36'd00000000;
					10'd0845: dataout<=36'd00000000;
					10'd0846: dataout<=36'd00000000;
					10'd0847: dataout<=36'd00000000;
					10'd0848: dataout<=36'd00000000;
					10'd0849: dataout<=36'd00000000;
					10'd0850: dataout<=36'd00000000;
					10'd0851: dataout<=36'd00000000;
					10'd0852: dataout<=36'd00000000;
					10'd0853: dataout<=36'd00000000;
					10'd0854: dataout<=36'd00000000;
					10'd0855: dataout<=36'd00000000;
					10'd0856: dataout<=36'd00000000;
					10'd0857: dataout<=36'd00000000;
					10'd0858: dataout<=36'd00000000;
					10'd0859: dataout<=36'd00000000;
					10'd0860: dataout<=36'd00000000;
					10'd0861: dataout<=36'd00000000;
					10'd0862: dataout<=36'd00000000;
					10'd0863: dataout<=36'd00000000;
					10'd0864: dataout<=36'd00000000;
					10'd0865: dataout<=36'd00000000;
					10'd0866: dataout<=36'd00000000;
					10'd0867: dataout<=36'd00000000;
					10'd0868: dataout<=36'd00000000;
					10'd0869: dataout<=36'd00000000;
					10'd0870: dataout<=36'd00000000;
					10'd0871: dataout<=36'd00000000;
					10'd0872: dataout<=36'd00000000;
					10'd0873: dataout<=36'd00000000;
					10'd0874: dataout<=36'd00000000;
					10'd0875: dataout<=36'd00000000;
					10'd0876: dataout<=36'd00000000;
					10'd0877: dataout<=36'd00000000;
					10'd0878: dataout<=36'd00000000;
					10'd0879: dataout<=36'd00000000;
					10'd0880: dataout<=36'd00000000;
					10'd0881: dataout<=36'd00000000;
					10'd0882: dataout<=36'd00000000;
					10'd0883: dataout<=36'd00000000;
					10'd0884: dataout<=36'd00000000;
					10'd0885: dataout<=36'd00000000;
					10'd0886: dataout<=36'd00000000;
					10'd0887: dataout<=36'd00000000;
					10'd0888: dataout<=36'd00000000;
					10'd0889: dataout<=36'd00000000;
					10'd0890: dataout<=36'd00000000;
					10'd0891: dataout<=36'd00000000;
					10'd0892: dataout<=36'd00000000;
					10'd0893: dataout<=36'd00000000;
					10'd0894: dataout<=36'd00000000;
					10'd0895: dataout<=36'd00000000;
					10'd0896: dataout<=36'd00000000;
					10'd0897: dataout<=36'd00000000;
					10'd0898: dataout<=36'd00000000;
					10'd0899: dataout<=36'd00000000;
					10'd0900: dataout<=36'd00000000;
					10'd0901: dataout<=36'd00000000;
					10'd0902: dataout<=36'd00000000;
					10'd0903: dataout<=36'd00000000;
					10'd0904: dataout<=36'd00000000;
					10'd0905: dataout<=36'd00000000;
					10'd0906: dataout<=36'd00000000;
					10'd0907: dataout<=36'd00000000;
					10'd0908: dataout<=36'd00000000;
					10'd0909: dataout<=36'd00000000;
					10'd0910: dataout<=36'd00000000;
					10'd0911: dataout<=36'd00000000;
					10'd0912: dataout<=36'd00000000;
					10'd0913: dataout<=36'd00000000;
					10'd0914: dataout<=36'd00000000;
					10'd0915: dataout<=36'd00000000;
					10'd0916: dataout<=36'd00000000;
					10'd0917: dataout<=36'd00000000;
					10'd0918: dataout<=36'd00000000;
					10'd0919: dataout<=36'd00000000;
					10'd0920: dataout<=36'd00000000;
					10'd0921: dataout<=36'd00000000;
					10'd0922: dataout<=36'd00000000;
					10'd0923: dataout<=36'd00000000;
					10'd0924: dataout<=36'd00000000;
					10'd0925: dataout<=36'd00000000;
					10'd0926: dataout<=36'd00000000;
					10'd0927: dataout<=36'd00000000;
					10'd0928: dataout<=36'd00000000;
					10'd0929: dataout<=36'd00000000;
					10'd0930: dataout<=36'd00000000;
					10'd0931: dataout<=36'd00000000;
					10'd0932: dataout<=36'd00000000;
					10'd0933: dataout<=36'd00000000;
					10'd0934: dataout<=36'd00000000;
					10'd0935: dataout<=36'd00000000;
					10'd0936: dataout<=36'd00000000;
					10'd0937: dataout<=36'd00000000;
					10'd0938: dataout<=36'd00000000;
					10'd0939: dataout<=36'd00000000;
					10'd0940: dataout<=36'd00000000;
					10'd0941: dataout<=36'd00000000;
					10'd0942: dataout<=36'd00000000;
					10'd0943: dataout<=36'd00000000;
					10'd0944: dataout<=36'd00000000;
					10'd0945: dataout<=36'd00000000;
					10'd0946: dataout<=36'd00000000;
					10'd0947: dataout<=36'd00000000;
					10'd0948: dataout<=36'd00000000;
					10'd0949: dataout<=36'd00000000;
					10'd0950: dataout<=36'd00000000;
					10'd0951: dataout<=36'd00000000;
					10'd0952: dataout<=36'd00000000;
					10'd0953: dataout<=36'd00000000;
					10'd0954: dataout<=36'd00000000;
					10'd0955: dataout<=36'd00000000;
					10'd0956: dataout<=36'd00000000;
					10'd0957: dataout<=36'd00000000;
					10'd0958: dataout<=36'd00000000;
					10'd0959: dataout<=36'd00000000;
					10'd0960: dataout<=36'd00000000;
					10'd0961: dataout<=36'd00000000;
					10'd0962: dataout<=36'd00000000;
					10'd0963: dataout<=36'd00000000;
					10'd0964: dataout<=36'd00000000;
					10'd0965: dataout<=36'd00000000;
					10'd0966: dataout<=36'd00000000;
					10'd0967: dataout<=36'd00000000;
					10'd0968: dataout<=36'd00000000;
					10'd0969: dataout<=36'd00000000;
					10'd0970: dataout<=36'd00000000;
					10'd0971: dataout<=36'd00000000;
					10'd0972: dataout<=36'd00000000;
					10'd0973: dataout<=36'd00000000;
					10'd0974: dataout<=36'd00000000;
					10'd0975: dataout<=36'd00000000;
					10'd0976: dataout<=36'd00000000;
					10'd0977: dataout<=36'd00000000;
					10'd0978: dataout<=36'd00000000;
					10'd0979: dataout<=36'd00000000;
					10'd0980: dataout<=36'd00000000;
					10'd0981: dataout<=36'd00000000;
					10'd0982: dataout<=36'd00000000;
					10'd0983: dataout<=36'd00000000;
					10'd0984: dataout<=36'd00000000;
					10'd0985: dataout<=36'd00000000;
					10'd0986: dataout<=36'd00000000;
					10'd0987: dataout<=36'd00000000;
					10'd0988: dataout<=36'd00000000;
					10'd0989: dataout<=36'd00000000;
					10'd0990: dataout<=36'd00000000;
					10'd0991: dataout<=36'd00000000;
					10'd0992: dataout<=36'd00000000;
					10'd0993: dataout<=36'd00000000;
					10'd0994: dataout<=36'd00000000;
					10'd0995: dataout<=36'd00000000;
					10'd0996: dataout<=36'd00000000;
					10'd0997: dataout<=36'd00000000;
					10'd0998: dataout<=36'd00000000;
					10'd0999: dataout<=36'd00000000;
					10'd1000: dataout<=36'd00000000;
					10'd1001: dataout<=36'd00000000;
					10'd1002: dataout<=36'd00000000;
					10'd1003: dataout<=36'd00000000;
					10'd1004: dataout<=36'd00000000;
					10'd1005: dataout<=36'd00000000;
					10'd1006: dataout<=36'd00000000;
					10'd1007: dataout<=36'd00000000;
					10'd1008: dataout<=36'd00000000;
					10'd1009: dataout<=36'd00000000;
					10'd1010: dataout<=36'd00000000;
					10'd1011: dataout<=36'd00000000;
					10'd1012: dataout<=36'd00000000;
					10'd1013: dataout<=36'd00000000;
					10'd1014: dataout<=36'd00000000;
					10'd1015: dataout<=36'd00000000;
					10'd1016: dataout<=36'd00000000;
					10'd1017: dataout<=36'd00000000;
					10'd1018: dataout<=36'd00000000;
					10'd1019: dataout<=36'd00000000;
					10'd1020: dataout<=36'd00000000;
					10'd1021: dataout<=36'd00000000;
					10'd1022: dataout<=36'd00000000;
					10'd1023: dataout<=36'd00000000;
				endcase
			end
		end
	end
endmodule

